
`include "nodeadder.v"

module LFPrefixSum128 (  // Ladner-Fischer
    input [127:0] mask,

    output [1023:0] psum
);

// Stage 1
wire [1:0] st1 [0:127];

assign st1[0]  = {1'b0, mask[0]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa1 (.a(mask[0]), .b(mask[1]), .y(st1[1]));
assign st1[2]  = {1'b0, mask[2]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa3 (.a(mask[2]), .b(mask[3]), .y(st1[3]));
assign st1[4]  = {1'b0, mask[4]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa5 (.a(mask[4]), .b(mask[5]), .y(st1[5]));
assign st1[6]  = {1'b0, mask[6]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa7 (.a(mask[6]), .b(mask[7]), .y(st1[7]));
assign st1[8]  = {1'b0, mask[8]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa9 (.a(mask[8]), .b(mask[9]), .y(st1[9]));
assign st1[10]  = {1'b0, mask[10]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa11 (.a(mask[10]), .b(mask[11]), .y(st1[11]));
assign st1[12]  = {1'b0, mask[12]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa13 (.a(mask[12]), .b(mask[13]), .y(st1[13]));
assign st1[14]  = {1'b0, mask[14]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa15 (.a(mask[14]), .b(mask[15]), .y(st1[15]));
assign st1[16]  = {1'b0, mask[16]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa17 (.a(mask[16]), .b(mask[17]), .y(st1[17]));
assign st1[18]  = {1'b0, mask[18]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa19 (.a(mask[18]), .b(mask[19]), .y(st1[19]));
assign st1[20]  = {1'b0, mask[20]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa21 (.a(mask[20]), .b(mask[21]), .y(st1[21]));
assign st1[22]  = {1'b0, mask[22]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa23 (.a(mask[22]), .b(mask[23]), .y(st1[23]));
assign st1[24]  = {1'b0, mask[24]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa25 (.a(mask[24]), .b(mask[25]), .y(st1[25]));
assign st1[26]  = {1'b0, mask[26]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa27 (.a(mask[26]), .b(mask[27]), .y(st1[27]));
assign st1[28]  = {1'b0, mask[28]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa29 (.a(mask[28]), .b(mask[29]), .y(st1[29]));
assign st1[30]  = {1'b0, mask[30]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa31 (.a(mask[30]), .b(mask[31]), .y(st1[31]));
assign st1[32]  = {1'b0, mask[32]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa33 (.a(mask[32]), .b(mask[33]), .y(st1[33]));
assign st1[34]  = {1'b0, mask[34]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa35 (.a(mask[34]), .b(mask[35]), .y(st1[35]));
assign st1[36]  = {1'b0, mask[36]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa37 (.a(mask[36]), .b(mask[37]), .y(st1[37]));
assign st1[38]  = {1'b0, mask[38]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa39 (.a(mask[38]), .b(mask[39]), .y(st1[39]));
assign st1[40]  = {1'b0, mask[40]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa41 (.a(mask[40]), .b(mask[41]), .y(st1[41]));
assign st1[42]  = {1'b0, mask[42]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa43 (.a(mask[42]), .b(mask[43]), .y(st1[43]));
assign st1[44]  = {1'b0, mask[44]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa45 (.a(mask[44]), .b(mask[45]), .y(st1[45]));
assign st1[46]  = {1'b0, mask[46]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa47 (.a(mask[46]), .b(mask[47]), .y(st1[47]));
assign st1[48]  = {1'b0, mask[48]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa49 (.a(mask[48]), .b(mask[49]), .y(st1[49]));
assign st1[50]  = {1'b0, mask[50]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa51 (.a(mask[50]), .b(mask[51]), .y(st1[51]));
assign st1[52]  = {1'b0, mask[52]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa53 (.a(mask[52]), .b(mask[53]), .y(st1[53]));
assign st1[54]  = {1'b0, mask[54]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa55 (.a(mask[54]), .b(mask[55]), .y(st1[55]));
assign st1[56]  = {1'b0, mask[56]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa57 (.a(mask[56]), .b(mask[57]), .y(st1[57]));
assign st1[58]  = {1'b0, mask[58]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa59 (.a(mask[58]), .b(mask[59]), .y(st1[59]));
assign st1[60]  = {1'b0, mask[60]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa61 (.a(mask[60]), .b(mask[61]), .y(st1[61]));
assign st1[62]  = {1'b0, mask[62]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa63 (.a(mask[62]), .b(mask[63]), .y(st1[63]));
assign st1[64]  = {1'b0, mask[64]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa65 (.a(mask[64]), .b(mask[65]), .y(st1[65]));
assign st1[66]  = {1'b0, mask[66]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa67 (.a(mask[66]), .b(mask[67]), .y(st1[67]));
assign st1[68]  = {1'b0, mask[68]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa69 (.a(mask[68]), .b(mask[69]), .y(st1[69]));
assign st1[70]  = {1'b0, mask[70]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa71 (.a(mask[70]), .b(mask[71]), .y(st1[71]));
assign st1[72]  = {1'b0, mask[72]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa73 (.a(mask[72]), .b(mask[73]), .y(st1[73]));
assign st1[74]  = {1'b0, mask[74]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa75 (.a(mask[74]), .b(mask[75]), .y(st1[75]));
assign st1[76]  = {1'b0, mask[76]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa77 (.a(mask[76]), .b(mask[77]), .y(st1[77]));
assign st1[78]  = {1'b0, mask[78]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa79 (.a(mask[78]), .b(mask[79]), .y(st1[79]));
assign st1[80]  = {1'b0, mask[80]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa81 (.a(mask[80]), .b(mask[81]), .y(st1[81]));
assign st1[82]  = {1'b0, mask[82]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa83 (.a(mask[82]), .b(mask[83]), .y(st1[83]));
assign st1[84]  = {1'b0, mask[84]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa85 (.a(mask[84]), .b(mask[85]), .y(st1[85]));
assign st1[86]  = {1'b0, mask[86]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa87 (.a(mask[86]), .b(mask[87]), .y(st1[87]));
assign st1[88]  = {1'b0, mask[88]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa89 (.a(mask[88]), .b(mask[89]), .y(st1[89]));
assign st1[90]  = {1'b0, mask[90]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa91 (.a(mask[90]), .b(mask[91]), .y(st1[91]));
assign st1[92]  = {1'b0, mask[92]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa93 (.a(mask[92]), .b(mask[93]), .y(st1[93]));
assign st1[94]  = {1'b0, mask[94]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa95 (.a(mask[94]), .b(mask[95]), .y(st1[95]));
assign st1[96]  = {1'b0, mask[96]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa97 (.a(mask[96]), .b(mask[97]), .y(st1[97]));
assign st1[98]  = {1'b0, mask[98]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa99 (.a(mask[98]), .b(mask[99]), .y(st1[99]));
assign st1[100]  = {1'b0, mask[100]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa101 (.a(mask[100]), .b(mask[101]), .y(st1[101]));
assign st1[102]  = {1'b0, mask[102]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa103 (.a(mask[102]), .b(mask[103]), .y(st1[103]));
assign st1[104]  = {1'b0, mask[104]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa105 (.a(mask[104]), .b(mask[105]), .y(st1[105]));
assign st1[106]  = {1'b0, mask[106]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa107 (.a(mask[106]), .b(mask[107]), .y(st1[107]));
assign st1[108]  = {1'b0, mask[108]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa109 (.a(mask[108]), .b(mask[109]), .y(st1[109]));
assign st1[110]  = {1'b0, mask[110]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa111 (.a(mask[110]), .b(mask[111]), .y(st1[111]));
assign st1[112]  = {1'b0, mask[112]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa113 (.a(mask[112]), .b(mask[113]), .y(st1[113]));
assign st1[114]  = {1'b0, mask[114]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa115 (.a(mask[114]), .b(mask[115]), .y(st1[115]));
assign st1[116]  = {1'b0, mask[116]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa117 (.a(mask[116]), .b(mask[117]), .y(st1[117]));
assign st1[118]  = {1'b0, mask[118]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa119 (.a(mask[118]), .b(mask[119]), .y(st1[119]));
assign st1[120]  = {1'b0, mask[120]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa121 (.a(mask[120]), .b(mask[121]), .y(st1[121]));
assign st1[122]  = {1'b0, mask[122]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa123 (.a(mask[122]), .b(mask[123]), .y(st1[123]));
assign st1[124]  = {1'b0, mask[124]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa125 (.a(mask[124]), .b(mask[125]), .y(st1[125]));
assign st1[126]  = {1'b0, mask[126]};
NodeAdder #(.WORD_WIDTH(1)) st1_pa127 (.a(mask[126]), .b(mask[127]), .y(st1[127]));



// Stage 2
wire [2:0] st2 [0:127];

assign st2[0]  = {1'b0, st1[0]};
assign st2[1]  = {1'b0, st1[1]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa2 (.a(st1[1]), .b(st1[2]), .y(st2[2]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa3 (.a(st1[1]), .b(st1[3]), .y(st2[3]));
assign st2[4]  = {1'b0, st1[4]};
assign st2[5]  = {1'b0, st1[5]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa6 (.a(st1[5]), .b(st1[6]), .y(st2[6]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa7 (.a(st1[5]), .b(st1[7]), .y(st2[7]));
assign st2[8]  = {1'b0, st1[8]};
assign st2[9]  = {1'b0, st1[9]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa10 (.a(st1[9]), .b(st1[10]), .y(st2[10]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa11 (.a(st1[9]), .b(st1[11]), .y(st2[11]));
assign st2[12]  = {1'b0, st1[12]};
assign st2[13]  = {1'b0, st1[13]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa14 (.a(st1[13]), .b(st1[14]), .y(st2[14]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa15 (.a(st1[13]), .b(st1[15]), .y(st2[15]));
assign st2[16]  = {1'b0, st1[16]};
assign st2[17]  = {1'b0, st1[17]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa18 (.a(st1[17]), .b(st1[18]), .y(st2[18]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa19 (.a(st1[17]), .b(st1[19]), .y(st2[19]));
assign st2[20]  = {1'b0, st1[20]};
assign st2[21]  = {1'b0, st1[21]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa22 (.a(st1[21]), .b(st1[22]), .y(st2[22]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa23 (.a(st1[21]), .b(st1[23]), .y(st2[23]));
assign st2[24]  = {1'b0, st1[24]};
assign st2[25]  = {1'b0, st1[25]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa26 (.a(st1[25]), .b(st1[26]), .y(st2[26]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa27 (.a(st1[25]), .b(st1[27]), .y(st2[27]));
assign st2[28]  = {1'b0, st1[28]};
assign st2[29]  = {1'b0, st1[29]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa30 (.a(st1[29]), .b(st1[30]), .y(st2[30]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa31 (.a(st1[29]), .b(st1[31]), .y(st2[31]));
assign st2[32]  = {1'b0, st1[32]};
assign st2[33]  = {1'b0, st1[33]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa34 (.a(st1[33]), .b(st1[34]), .y(st2[34]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa35 (.a(st1[33]), .b(st1[35]), .y(st2[35]));
assign st2[36]  = {1'b0, st1[36]};
assign st2[37]  = {1'b0, st1[37]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa38 (.a(st1[37]), .b(st1[38]), .y(st2[38]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa39 (.a(st1[37]), .b(st1[39]), .y(st2[39]));
assign st2[40]  = {1'b0, st1[40]};
assign st2[41]  = {1'b0, st1[41]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa42 (.a(st1[41]), .b(st1[42]), .y(st2[42]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa43 (.a(st1[41]), .b(st1[43]), .y(st2[43]));
assign st2[44]  = {1'b0, st1[44]};
assign st2[45]  = {1'b0, st1[45]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa46 (.a(st1[45]), .b(st1[46]), .y(st2[46]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa47 (.a(st1[45]), .b(st1[47]), .y(st2[47]));
assign st2[48]  = {1'b0, st1[48]};
assign st2[49]  = {1'b0, st1[49]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa50 (.a(st1[49]), .b(st1[50]), .y(st2[50]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa51 (.a(st1[49]), .b(st1[51]), .y(st2[51]));
assign st2[52]  = {1'b0, st1[52]};
assign st2[53]  = {1'b0, st1[53]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa54 (.a(st1[53]), .b(st1[54]), .y(st2[54]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa55 (.a(st1[53]), .b(st1[55]), .y(st2[55]));
assign st2[56]  = {1'b0, st1[56]};
assign st2[57]  = {1'b0, st1[57]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa58 (.a(st1[57]), .b(st1[58]), .y(st2[58]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa59 (.a(st1[57]), .b(st1[59]), .y(st2[59]));
assign st2[60]  = {1'b0, st1[60]};
assign st2[61]  = {1'b0, st1[61]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa62 (.a(st1[61]), .b(st1[62]), .y(st2[62]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa63 (.a(st1[61]), .b(st1[63]), .y(st2[63]));
assign st2[64]  = {1'b0, st1[64]};
assign st2[65]  = {1'b0, st1[65]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa66 (.a(st1[65]), .b(st1[66]), .y(st2[66]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa67 (.a(st1[65]), .b(st1[67]), .y(st2[67]));
assign st2[68]  = {1'b0, st1[68]};
assign st2[69]  = {1'b0, st1[69]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa70 (.a(st1[69]), .b(st1[70]), .y(st2[70]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa71 (.a(st1[69]), .b(st1[71]), .y(st2[71]));
assign st2[72]  = {1'b0, st1[72]};
assign st2[73]  = {1'b0, st1[73]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa74 (.a(st1[73]), .b(st1[74]), .y(st2[74]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa75 (.a(st1[73]), .b(st1[75]), .y(st2[75]));
assign st2[76]  = {1'b0, st1[76]};
assign st2[77]  = {1'b0, st1[77]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa78 (.a(st1[77]), .b(st1[78]), .y(st2[78]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa79 (.a(st1[77]), .b(st1[79]), .y(st2[79]));
assign st2[80]  = {1'b0, st1[80]};
assign st2[81]  = {1'b0, st1[81]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa82 (.a(st1[81]), .b(st1[82]), .y(st2[82]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa83 (.a(st1[81]), .b(st1[83]), .y(st2[83]));
assign st2[84]  = {1'b0, st1[84]};
assign st2[85]  = {1'b0, st1[85]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa86 (.a(st1[85]), .b(st1[86]), .y(st2[86]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa87 (.a(st1[85]), .b(st1[87]), .y(st2[87]));
assign st2[88]  = {1'b0, st1[88]};
assign st2[89]  = {1'b0, st1[89]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa90 (.a(st1[89]), .b(st1[90]), .y(st2[90]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa91 (.a(st1[89]), .b(st1[91]), .y(st2[91]));
assign st2[92]  = {1'b0, st1[92]};
assign st2[93]  = {1'b0, st1[93]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa94 (.a(st1[93]), .b(st1[94]), .y(st2[94]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa95 (.a(st1[93]), .b(st1[95]), .y(st2[95]));
assign st2[96]  = {1'b0, st1[96]};
assign st2[97]  = {1'b0, st1[97]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa98 (.a(st1[97]), .b(st1[98]), .y(st2[98]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa99 (.a(st1[97]), .b(st1[99]), .y(st2[99]));
assign st2[100]  = {1'b0, st1[100]};
assign st2[101]  = {1'b0, st1[101]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa102 (.a(st1[101]), .b(st1[102]), .y(st2[102]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa103 (.a(st1[101]), .b(st1[103]), .y(st2[103]));
assign st2[104]  = {1'b0, st1[104]};
assign st2[105]  = {1'b0, st1[105]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa106 (.a(st1[105]), .b(st1[106]), .y(st2[106]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa107 (.a(st1[105]), .b(st1[107]), .y(st2[107]));
assign st2[108]  = {1'b0, st1[108]};
assign st2[109]  = {1'b0, st1[109]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa110 (.a(st1[109]), .b(st1[110]), .y(st2[110]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa111 (.a(st1[109]), .b(st1[111]), .y(st2[111]));
assign st2[112]  = {1'b0, st1[112]};
assign st2[113]  = {1'b0, st1[113]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa114 (.a(st1[113]), .b(st1[114]), .y(st2[114]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa115 (.a(st1[113]), .b(st1[115]), .y(st2[115]));
assign st2[116]  = {1'b0, st1[116]};
assign st2[117]  = {1'b0, st1[117]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa118 (.a(st1[117]), .b(st1[118]), .y(st2[118]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa119 (.a(st1[117]), .b(st1[119]), .y(st2[119]));
assign st2[120]  = {1'b0, st1[120]};
assign st2[121]  = {1'b0, st1[121]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa122 (.a(st1[121]), .b(st1[122]), .y(st2[122]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa123 (.a(st1[121]), .b(st1[123]), .y(st2[123]));
assign st2[124]  = {1'b0, st1[124]};
assign st2[125]  = {1'b0, st1[125]};
NodeAdder #(.WORD_WIDTH(2)) st2_pa126 (.a(st1[125]), .b(st1[126]), .y(st2[126]));
NodeAdder #(.WORD_WIDTH(2)) st2_pa127 (.a(st1[125]), .b(st1[127]), .y(st2[127]));



// Stage 3
wire [3:0] st3 [0:127];

assign st3[0]  = {1'b0, st2[0]};
assign st3[1]  = {1'b0, st2[1]};
assign st3[2]  = {1'b0, st2[2]};
assign st3[3]  = {1'b0, st2[3]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa4 (.a(st2[3]), .b(st2[4]), .y(st3[4]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa5 (.a(st2[3]), .b(st2[5]), .y(st3[5]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa6 (.a(st2[3]), .b(st2[6]), .y(st3[6]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa7 (.a(st2[3]), .b(st2[7]), .y(st3[7]));
assign st3[8]  = {1'b0, st2[8]};
assign st3[9]  = {1'b0, st2[9]};
assign st3[10]  = {1'b0, st2[10]};
assign st3[11]  = {1'b0, st2[11]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa12 (.a(st2[11]), .b(st2[12]), .y(st3[12]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa13 (.a(st2[11]), .b(st2[13]), .y(st3[13]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa14 (.a(st2[11]), .b(st2[14]), .y(st3[14]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa15 (.a(st2[11]), .b(st2[15]), .y(st3[15]));
assign st3[16]  = {1'b0, st2[16]};
assign st3[17]  = {1'b0, st2[17]};
assign st3[18]  = {1'b0, st2[18]};
assign st3[19]  = {1'b0, st2[19]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa20 (.a(st2[19]), .b(st2[20]), .y(st3[20]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa21 (.a(st2[19]), .b(st2[21]), .y(st3[21]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa22 (.a(st2[19]), .b(st2[22]), .y(st3[22]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa23 (.a(st2[19]), .b(st2[23]), .y(st3[23]));
assign st3[24]  = {1'b0, st2[24]};
assign st3[25]  = {1'b0, st2[25]};
assign st3[26]  = {1'b0, st2[26]};
assign st3[27]  = {1'b0, st2[27]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa28 (.a(st2[27]), .b(st2[28]), .y(st3[28]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa29 (.a(st2[27]), .b(st2[29]), .y(st3[29]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa30 (.a(st2[27]), .b(st2[30]), .y(st3[30]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa31 (.a(st2[27]), .b(st2[31]), .y(st3[31]));
assign st3[32]  = {1'b0, st2[32]};
assign st3[33]  = {1'b0, st2[33]};
assign st3[34]  = {1'b0, st2[34]};
assign st3[35]  = {1'b0, st2[35]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa36 (.a(st2[35]), .b(st2[36]), .y(st3[36]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa37 (.a(st2[35]), .b(st2[37]), .y(st3[37]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa38 (.a(st2[35]), .b(st2[38]), .y(st3[38]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa39 (.a(st2[35]), .b(st2[39]), .y(st3[39]));
assign st3[40]  = {1'b0, st2[40]};
assign st3[41]  = {1'b0, st2[41]};
assign st3[42]  = {1'b0, st2[42]};
assign st3[43]  = {1'b0, st2[43]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa44 (.a(st2[43]), .b(st2[44]), .y(st3[44]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa45 (.a(st2[43]), .b(st2[45]), .y(st3[45]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa46 (.a(st2[43]), .b(st2[46]), .y(st3[46]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa47 (.a(st2[43]), .b(st2[47]), .y(st3[47]));
assign st3[48]  = {1'b0, st2[48]};
assign st3[49]  = {1'b0, st2[49]};
assign st3[50]  = {1'b0, st2[50]};
assign st3[51]  = {1'b0, st2[51]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa52 (.a(st2[51]), .b(st2[52]), .y(st3[52]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa53 (.a(st2[51]), .b(st2[53]), .y(st3[53]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa54 (.a(st2[51]), .b(st2[54]), .y(st3[54]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa55 (.a(st2[51]), .b(st2[55]), .y(st3[55]));
assign st3[56]  = {1'b0, st2[56]};
assign st3[57]  = {1'b0, st2[57]};
assign st3[58]  = {1'b0, st2[58]};
assign st3[59]  = {1'b0, st2[59]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa60 (.a(st2[59]), .b(st2[60]), .y(st3[60]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa61 (.a(st2[59]), .b(st2[61]), .y(st3[61]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa62 (.a(st2[59]), .b(st2[62]), .y(st3[62]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa63 (.a(st2[59]), .b(st2[63]), .y(st3[63]));
assign st3[64]  = {1'b0, st2[64]};
assign st3[65]  = {1'b0, st2[65]};
assign st3[66]  = {1'b0, st2[66]};
assign st3[67]  = {1'b0, st2[67]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa68 (.a(st2[67]), .b(st2[68]), .y(st3[68]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa69 (.a(st2[67]), .b(st2[69]), .y(st3[69]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa70 (.a(st2[67]), .b(st2[70]), .y(st3[70]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa71 (.a(st2[67]), .b(st2[71]), .y(st3[71]));
assign st3[72]  = {1'b0, st2[72]};
assign st3[73]  = {1'b0, st2[73]};
assign st3[74]  = {1'b0, st2[74]};
assign st3[75]  = {1'b0, st2[75]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa76 (.a(st2[75]), .b(st2[76]), .y(st3[76]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa77 (.a(st2[75]), .b(st2[77]), .y(st3[77]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa78 (.a(st2[75]), .b(st2[78]), .y(st3[78]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa79 (.a(st2[75]), .b(st2[79]), .y(st3[79]));
assign st3[80]  = {1'b0, st2[80]};
assign st3[81]  = {1'b0, st2[81]};
assign st3[82]  = {1'b0, st2[82]};
assign st3[83]  = {1'b0, st2[83]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa84 (.a(st2[83]), .b(st2[84]), .y(st3[84]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa85 (.a(st2[83]), .b(st2[85]), .y(st3[85]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa86 (.a(st2[83]), .b(st2[86]), .y(st3[86]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa87 (.a(st2[83]), .b(st2[87]), .y(st3[87]));
assign st3[88]  = {1'b0, st2[88]};
assign st3[89]  = {1'b0, st2[89]};
assign st3[90]  = {1'b0, st2[90]};
assign st3[91]  = {1'b0, st2[91]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa92 (.a(st2[91]), .b(st2[92]), .y(st3[92]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa93 (.a(st2[91]), .b(st2[93]), .y(st3[93]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa94 (.a(st2[91]), .b(st2[94]), .y(st3[94]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa95 (.a(st2[91]), .b(st2[95]), .y(st3[95]));
assign st3[96]  = {1'b0, st2[96]};
assign st3[97]  = {1'b0, st2[97]};
assign st3[98]  = {1'b0, st2[98]};
assign st3[99]  = {1'b0, st2[99]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa100 (.a(st2[99]), .b(st2[100]), .y(st3[100]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa101 (.a(st2[99]), .b(st2[101]), .y(st3[101]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa102 (.a(st2[99]), .b(st2[102]), .y(st3[102]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa103 (.a(st2[99]), .b(st2[103]), .y(st3[103]));
assign st3[104]  = {1'b0, st2[104]};
assign st3[105]  = {1'b0, st2[105]};
assign st3[106]  = {1'b0, st2[106]};
assign st3[107]  = {1'b0, st2[107]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa108 (.a(st2[107]), .b(st2[108]), .y(st3[108]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa109 (.a(st2[107]), .b(st2[109]), .y(st3[109]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa110 (.a(st2[107]), .b(st2[110]), .y(st3[110]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa111 (.a(st2[107]), .b(st2[111]), .y(st3[111]));
assign st3[112]  = {1'b0, st2[112]};
assign st3[113]  = {1'b0, st2[113]};
assign st3[114]  = {1'b0, st2[114]};
assign st3[115]  = {1'b0, st2[115]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa116 (.a(st2[115]), .b(st2[116]), .y(st3[116]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa117 (.a(st2[115]), .b(st2[117]), .y(st3[117]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa118 (.a(st2[115]), .b(st2[118]), .y(st3[118]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa119 (.a(st2[115]), .b(st2[119]), .y(st3[119]));
assign st3[120]  = {1'b0, st2[120]};
assign st3[121]  = {1'b0, st2[121]};
assign st3[122]  = {1'b0, st2[122]};
assign st3[123]  = {1'b0, st2[123]};
NodeAdder #(.WORD_WIDTH(3)) st3_pa124 (.a(st2[123]), .b(st2[124]), .y(st3[124]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa125 (.a(st2[123]), .b(st2[125]), .y(st3[125]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa126 (.a(st2[123]), .b(st2[126]), .y(st3[126]));
NodeAdder #(.WORD_WIDTH(3)) st3_pa127 (.a(st2[123]), .b(st2[127]), .y(st3[127]));



// Stage 4
wire [4:0] st4 [0:127];

assign st4[0]  = {1'b0, st3[0]};
assign st4[1]  = {1'b0, st3[1]};
assign st4[2]  = {1'b0, st3[2]};
assign st4[3]  = {1'b0, st3[3]};
assign st4[4]  = {1'b0, st3[4]};
assign st4[5]  = {1'b0, st3[5]};
assign st4[6]  = {1'b0, st3[6]};
assign st4[7]  = {1'b0, st3[7]};
NodeAdder #(.WORD_WIDTH(4)) st4_pa8 (.a(st3[7]), .b(st3[8]), .y(st4[8]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa9 (.a(st3[7]), .b(st3[9]), .y(st4[9]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa10 (.a(st3[7]), .b(st3[10]), .y(st4[10]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa11 (.a(st3[7]), .b(st3[11]), .y(st4[11]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa12 (.a(st3[7]), .b(st3[12]), .y(st4[12]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa13 (.a(st3[7]), .b(st3[13]), .y(st4[13]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa14 (.a(st3[7]), .b(st3[14]), .y(st4[14]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa15 (.a(st3[7]), .b(st3[15]), .y(st4[15]));
assign st4[16]  = {1'b0, st3[16]};
assign st4[17]  = {1'b0, st3[17]};
assign st4[18]  = {1'b0, st3[18]};
assign st4[19]  = {1'b0, st3[19]};
assign st4[20]  = {1'b0, st3[20]};
assign st4[21]  = {1'b0, st3[21]};
assign st4[22]  = {1'b0, st3[22]};
assign st4[23]  = {1'b0, st3[23]};
NodeAdder #(.WORD_WIDTH(4)) st4_pa24 (.a(st3[23]), .b(st3[24]), .y(st4[24]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa25 (.a(st3[23]), .b(st3[25]), .y(st4[25]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa26 (.a(st3[23]), .b(st3[26]), .y(st4[26]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa27 (.a(st3[23]), .b(st3[27]), .y(st4[27]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa28 (.a(st3[23]), .b(st3[28]), .y(st4[28]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa29 (.a(st3[23]), .b(st3[29]), .y(st4[29]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa30 (.a(st3[23]), .b(st3[30]), .y(st4[30]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa31 (.a(st3[23]), .b(st3[31]), .y(st4[31]));
assign st4[32]  = {1'b0, st3[32]};
assign st4[33]  = {1'b0, st3[33]};
assign st4[34]  = {1'b0, st3[34]};
assign st4[35]  = {1'b0, st3[35]};
assign st4[36]  = {1'b0, st3[36]};
assign st4[37]  = {1'b0, st3[37]};
assign st4[38]  = {1'b0, st3[38]};
assign st4[39]  = {1'b0, st3[39]};
NodeAdder #(.WORD_WIDTH(4)) st4_pa40 (.a(st3[39]), .b(st3[40]), .y(st4[40]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa41 (.a(st3[39]), .b(st3[41]), .y(st4[41]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa42 (.a(st3[39]), .b(st3[42]), .y(st4[42]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa43 (.a(st3[39]), .b(st3[43]), .y(st4[43]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa44 (.a(st3[39]), .b(st3[44]), .y(st4[44]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa45 (.a(st3[39]), .b(st3[45]), .y(st4[45]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa46 (.a(st3[39]), .b(st3[46]), .y(st4[46]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa47 (.a(st3[39]), .b(st3[47]), .y(st4[47]));
assign st4[48]  = {1'b0, st3[48]};
assign st4[49]  = {1'b0, st3[49]};
assign st4[50]  = {1'b0, st3[50]};
assign st4[51]  = {1'b0, st3[51]};
assign st4[52]  = {1'b0, st3[52]};
assign st4[53]  = {1'b0, st3[53]};
assign st4[54]  = {1'b0, st3[54]};
assign st4[55]  = {1'b0, st3[55]};
NodeAdder #(.WORD_WIDTH(4)) st4_pa56 (.a(st3[55]), .b(st3[56]), .y(st4[56]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa57 (.a(st3[55]), .b(st3[57]), .y(st4[57]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa58 (.a(st3[55]), .b(st3[58]), .y(st4[58]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa59 (.a(st3[55]), .b(st3[59]), .y(st4[59]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa60 (.a(st3[55]), .b(st3[60]), .y(st4[60]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa61 (.a(st3[55]), .b(st3[61]), .y(st4[61]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa62 (.a(st3[55]), .b(st3[62]), .y(st4[62]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa63 (.a(st3[55]), .b(st3[63]), .y(st4[63]));
assign st4[64]  = {1'b0, st3[64]};
assign st4[65]  = {1'b0, st3[65]};
assign st4[66]  = {1'b0, st3[66]};
assign st4[67]  = {1'b0, st3[67]};
assign st4[68]  = {1'b0, st3[68]};
assign st4[69]  = {1'b0, st3[69]};
assign st4[70]  = {1'b0, st3[70]};
assign st4[71]  = {1'b0, st3[71]};
NodeAdder #(.WORD_WIDTH(4)) st4_pa72 (.a(st3[71]), .b(st3[72]), .y(st4[72]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa73 (.a(st3[71]), .b(st3[73]), .y(st4[73]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa74 (.a(st3[71]), .b(st3[74]), .y(st4[74]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa75 (.a(st3[71]), .b(st3[75]), .y(st4[75]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa76 (.a(st3[71]), .b(st3[76]), .y(st4[76]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa77 (.a(st3[71]), .b(st3[77]), .y(st4[77]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa78 (.a(st3[71]), .b(st3[78]), .y(st4[78]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa79 (.a(st3[71]), .b(st3[79]), .y(st4[79]));
assign st4[80]  = {1'b0, st3[80]};
assign st4[81]  = {1'b0, st3[81]};
assign st4[82]  = {1'b0, st3[82]};
assign st4[83]  = {1'b0, st3[83]};
assign st4[84]  = {1'b0, st3[84]};
assign st4[85]  = {1'b0, st3[85]};
assign st4[86]  = {1'b0, st3[86]};
assign st4[87]  = {1'b0, st3[87]};
NodeAdder #(.WORD_WIDTH(4)) st4_pa88 (.a(st3[87]), .b(st3[88]), .y(st4[88]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa89 (.a(st3[87]), .b(st3[89]), .y(st4[89]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa90 (.a(st3[87]), .b(st3[90]), .y(st4[90]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa91 (.a(st3[87]), .b(st3[91]), .y(st4[91]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa92 (.a(st3[87]), .b(st3[92]), .y(st4[92]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa93 (.a(st3[87]), .b(st3[93]), .y(st4[93]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa94 (.a(st3[87]), .b(st3[94]), .y(st4[94]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa95 (.a(st3[87]), .b(st3[95]), .y(st4[95]));
assign st4[96]  = {1'b0, st3[96]};
assign st4[97]  = {1'b0, st3[97]};
assign st4[98]  = {1'b0, st3[98]};
assign st4[99]  = {1'b0, st3[99]};
assign st4[100]  = {1'b0, st3[100]};
assign st4[101]  = {1'b0, st3[101]};
assign st4[102]  = {1'b0, st3[102]};
assign st4[103]  = {1'b0, st3[103]};
NodeAdder #(.WORD_WIDTH(4)) st4_pa104 (.a(st3[103]), .b(st3[104]), .y(st4[104]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa105 (.a(st3[103]), .b(st3[105]), .y(st4[105]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa106 (.a(st3[103]), .b(st3[106]), .y(st4[106]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa107 (.a(st3[103]), .b(st3[107]), .y(st4[107]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa108 (.a(st3[103]), .b(st3[108]), .y(st4[108]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa109 (.a(st3[103]), .b(st3[109]), .y(st4[109]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa110 (.a(st3[103]), .b(st3[110]), .y(st4[110]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa111 (.a(st3[103]), .b(st3[111]), .y(st4[111]));
assign st4[112]  = {1'b0, st3[112]};
assign st4[113]  = {1'b0, st3[113]};
assign st4[114]  = {1'b0, st3[114]};
assign st4[115]  = {1'b0, st3[115]};
assign st4[116]  = {1'b0, st3[116]};
assign st4[117]  = {1'b0, st3[117]};
assign st4[118]  = {1'b0, st3[118]};
assign st4[119]  = {1'b0, st3[119]};
NodeAdder #(.WORD_WIDTH(4)) st4_pa120 (.a(st3[119]), .b(st3[120]), .y(st4[120]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa121 (.a(st3[119]), .b(st3[121]), .y(st4[121]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa122 (.a(st3[119]), .b(st3[122]), .y(st4[122]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa123 (.a(st3[119]), .b(st3[123]), .y(st4[123]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa124 (.a(st3[119]), .b(st3[124]), .y(st4[124]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa125 (.a(st3[119]), .b(st3[125]), .y(st4[125]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa126 (.a(st3[119]), .b(st3[126]), .y(st4[126]));
NodeAdder #(.WORD_WIDTH(4)) st4_pa127 (.a(st3[119]), .b(st3[127]), .y(st4[127]));



// Stage 5
wire [5:0] st5 [0:127];

assign st5[0]  = {1'b0, st4[0]};
assign st5[1]  = {1'b0, st4[1]};
assign st5[2]  = {1'b0, st4[2]};
assign st5[3]  = {1'b0, st4[3]};
assign st5[4]  = {1'b0, st4[4]};
assign st5[5]  = {1'b0, st4[5]};
assign st5[6]  = {1'b0, st4[6]};
assign st5[7]  = {1'b0, st4[7]};
assign st5[8]  = {1'b0, st4[8]};
assign st5[9]  = {1'b0, st4[9]};
assign st5[10]  = {1'b0, st4[10]};
assign st5[11]  = {1'b0, st4[11]};
assign st5[12]  = {1'b0, st4[12]};
assign st5[13]  = {1'b0, st4[13]};
assign st5[14]  = {1'b0, st4[14]};
assign st5[15]  = {1'b0, st4[15]};
NodeAdder #(.WORD_WIDTH(5)) st5_pa16 (.a(st4[15]), .b(st4[16]), .y(st5[16]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa17 (.a(st4[15]), .b(st4[17]), .y(st5[17]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa18 (.a(st4[15]), .b(st4[18]), .y(st5[18]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa19 (.a(st4[15]), .b(st4[19]), .y(st5[19]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa20 (.a(st4[15]), .b(st4[20]), .y(st5[20]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa21 (.a(st4[15]), .b(st4[21]), .y(st5[21]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa22 (.a(st4[15]), .b(st4[22]), .y(st5[22]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa23 (.a(st4[15]), .b(st4[23]), .y(st5[23]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa24 (.a(st4[15]), .b(st4[24]), .y(st5[24]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa25 (.a(st4[15]), .b(st4[25]), .y(st5[25]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa26 (.a(st4[15]), .b(st4[26]), .y(st5[26]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa27 (.a(st4[15]), .b(st4[27]), .y(st5[27]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa28 (.a(st4[15]), .b(st4[28]), .y(st5[28]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa29 (.a(st4[15]), .b(st4[29]), .y(st5[29]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa30 (.a(st4[15]), .b(st4[30]), .y(st5[30]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa31 (.a(st4[15]), .b(st4[31]), .y(st5[31]));
assign st5[32]  = {1'b0, st4[32]};
assign st5[33]  = {1'b0, st4[33]};
assign st5[34]  = {1'b0, st4[34]};
assign st5[35]  = {1'b0, st4[35]};
assign st5[36]  = {1'b0, st4[36]};
assign st5[37]  = {1'b0, st4[37]};
assign st5[38]  = {1'b0, st4[38]};
assign st5[39]  = {1'b0, st4[39]};
assign st5[40]  = {1'b0, st4[40]};
assign st5[41]  = {1'b0, st4[41]};
assign st5[42]  = {1'b0, st4[42]};
assign st5[43]  = {1'b0, st4[43]};
assign st5[44]  = {1'b0, st4[44]};
assign st5[45]  = {1'b0, st4[45]};
assign st5[46]  = {1'b0, st4[46]};
assign st5[47]  = {1'b0, st4[47]};
NodeAdder #(.WORD_WIDTH(5)) st5_pa48 (.a(st4[47]), .b(st4[48]), .y(st5[48]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa49 (.a(st4[47]), .b(st4[49]), .y(st5[49]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa50 (.a(st4[47]), .b(st4[50]), .y(st5[50]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa51 (.a(st4[47]), .b(st4[51]), .y(st5[51]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa52 (.a(st4[47]), .b(st4[52]), .y(st5[52]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa53 (.a(st4[47]), .b(st4[53]), .y(st5[53]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa54 (.a(st4[47]), .b(st4[54]), .y(st5[54]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa55 (.a(st4[47]), .b(st4[55]), .y(st5[55]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa56 (.a(st4[47]), .b(st4[56]), .y(st5[56]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa57 (.a(st4[47]), .b(st4[57]), .y(st5[57]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa58 (.a(st4[47]), .b(st4[58]), .y(st5[58]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa59 (.a(st4[47]), .b(st4[59]), .y(st5[59]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa60 (.a(st4[47]), .b(st4[60]), .y(st5[60]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa61 (.a(st4[47]), .b(st4[61]), .y(st5[61]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa62 (.a(st4[47]), .b(st4[62]), .y(st5[62]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa63 (.a(st4[47]), .b(st4[63]), .y(st5[63]));
assign st5[64]  = {1'b0, st4[64]};
assign st5[65]  = {1'b0, st4[65]};
assign st5[66]  = {1'b0, st4[66]};
assign st5[67]  = {1'b0, st4[67]};
assign st5[68]  = {1'b0, st4[68]};
assign st5[69]  = {1'b0, st4[69]};
assign st5[70]  = {1'b0, st4[70]};
assign st5[71]  = {1'b0, st4[71]};
assign st5[72]  = {1'b0, st4[72]};
assign st5[73]  = {1'b0, st4[73]};
assign st5[74]  = {1'b0, st4[74]};
assign st5[75]  = {1'b0, st4[75]};
assign st5[76]  = {1'b0, st4[76]};
assign st5[77]  = {1'b0, st4[77]};
assign st5[78]  = {1'b0, st4[78]};
assign st5[79]  = {1'b0, st4[79]};
NodeAdder #(.WORD_WIDTH(5)) st5_pa80 (.a(st4[79]), .b(st4[80]), .y(st5[80]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa81 (.a(st4[79]), .b(st4[81]), .y(st5[81]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa82 (.a(st4[79]), .b(st4[82]), .y(st5[82]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa83 (.a(st4[79]), .b(st4[83]), .y(st5[83]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa84 (.a(st4[79]), .b(st4[84]), .y(st5[84]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa85 (.a(st4[79]), .b(st4[85]), .y(st5[85]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa86 (.a(st4[79]), .b(st4[86]), .y(st5[86]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa87 (.a(st4[79]), .b(st4[87]), .y(st5[87]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa88 (.a(st4[79]), .b(st4[88]), .y(st5[88]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa89 (.a(st4[79]), .b(st4[89]), .y(st5[89]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa90 (.a(st4[79]), .b(st4[90]), .y(st5[90]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa91 (.a(st4[79]), .b(st4[91]), .y(st5[91]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa92 (.a(st4[79]), .b(st4[92]), .y(st5[92]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa93 (.a(st4[79]), .b(st4[93]), .y(st5[93]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa94 (.a(st4[79]), .b(st4[94]), .y(st5[94]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa95 (.a(st4[79]), .b(st4[95]), .y(st5[95]));
assign st5[96]  = {1'b0, st4[96]};
assign st5[97]  = {1'b0, st4[97]};
assign st5[98]  = {1'b0, st4[98]};
assign st5[99]  = {1'b0, st4[99]};
assign st5[100]  = {1'b0, st4[100]};
assign st5[101]  = {1'b0, st4[101]};
assign st5[102]  = {1'b0, st4[102]};
assign st5[103]  = {1'b0, st4[103]};
assign st5[104]  = {1'b0, st4[104]};
assign st5[105]  = {1'b0, st4[105]};
assign st5[106]  = {1'b0, st4[106]};
assign st5[107]  = {1'b0, st4[107]};
assign st5[108]  = {1'b0, st4[108]};
assign st5[109]  = {1'b0, st4[109]};
assign st5[110]  = {1'b0, st4[110]};
assign st5[111]  = {1'b0, st4[111]};
NodeAdder #(.WORD_WIDTH(5)) st5_pa112 (.a(st4[111]), .b(st4[112]), .y(st5[112]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa113 (.a(st4[111]), .b(st4[113]), .y(st5[113]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa114 (.a(st4[111]), .b(st4[114]), .y(st5[114]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa115 (.a(st4[111]), .b(st4[115]), .y(st5[115]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa116 (.a(st4[111]), .b(st4[116]), .y(st5[116]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa117 (.a(st4[111]), .b(st4[117]), .y(st5[117]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa118 (.a(st4[111]), .b(st4[118]), .y(st5[118]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa119 (.a(st4[111]), .b(st4[119]), .y(st5[119]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa120 (.a(st4[111]), .b(st4[120]), .y(st5[120]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa121 (.a(st4[111]), .b(st4[121]), .y(st5[121]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa122 (.a(st4[111]), .b(st4[122]), .y(st5[122]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa123 (.a(st4[111]), .b(st4[123]), .y(st5[123]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa124 (.a(st4[111]), .b(st4[124]), .y(st5[124]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa125 (.a(st4[111]), .b(st4[125]), .y(st5[125]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa126 (.a(st4[111]), .b(st4[126]), .y(st5[126]));
NodeAdder #(.WORD_WIDTH(5)) st5_pa127 (.a(st4[111]), .b(st4[127]), .y(st5[127]));



// Stage 6
wire [6:0] st6 [0:127];

assign st6[0]  = {1'b0, st5[0]};
assign st6[1]  = {1'b0, st5[1]};
assign st6[2]  = {1'b0, st5[2]};
assign st6[3]  = {1'b0, st5[3]};
assign st6[4]  = {1'b0, st5[4]};
assign st6[5]  = {1'b0, st5[5]};
assign st6[6]  = {1'b0, st5[6]};
assign st6[7]  = {1'b0, st5[7]};
assign st6[8]  = {1'b0, st5[8]};
assign st6[9]  = {1'b0, st5[9]};
assign st6[10]  = {1'b0, st5[10]};
assign st6[11]  = {1'b0, st5[11]};
assign st6[12]  = {1'b0, st5[12]};
assign st6[13]  = {1'b0, st5[13]};
assign st6[14]  = {1'b0, st5[14]};
assign st6[15]  = {1'b0, st5[15]};
assign st6[16]  = {1'b0, st5[16]};
assign st6[17]  = {1'b0, st5[17]};
assign st6[18]  = {1'b0, st5[18]};
assign st6[19]  = {1'b0, st5[19]};
assign st6[20]  = {1'b0, st5[20]};
assign st6[21]  = {1'b0, st5[21]};
assign st6[22]  = {1'b0, st5[22]};
assign st6[23]  = {1'b0, st5[23]};
assign st6[24]  = {1'b0, st5[24]};
assign st6[25]  = {1'b0, st5[25]};
assign st6[26]  = {1'b0, st5[26]};
assign st6[27]  = {1'b0, st5[27]};
assign st6[28]  = {1'b0, st5[28]};
assign st6[29]  = {1'b0, st5[29]};
assign st6[30]  = {1'b0, st5[30]};
assign st6[31]  = {1'b0, st5[31]};
NodeAdder #(.WORD_WIDTH(6)) st6_pa32 (.a(st5[31]), .b(st5[32]), .y(st6[32]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa33 (.a(st5[31]), .b(st5[33]), .y(st6[33]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa34 (.a(st5[31]), .b(st5[34]), .y(st6[34]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa35 (.a(st5[31]), .b(st5[35]), .y(st6[35]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa36 (.a(st5[31]), .b(st5[36]), .y(st6[36]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa37 (.a(st5[31]), .b(st5[37]), .y(st6[37]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa38 (.a(st5[31]), .b(st5[38]), .y(st6[38]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa39 (.a(st5[31]), .b(st5[39]), .y(st6[39]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa40 (.a(st5[31]), .b(st5[40]), .y(st6[40]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa41 (.a(st5[31]), .b(st5[41]), .y(st6[41]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa42 (.a(st5[31]), .b(st5[42]), .y(st6[42]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa43 (.a(st5[31]), .b(st5[43]), .y(st6[43]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa44 (.a(st5[31]), .b(st5[44]), .y(st6[44]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa45 (.a(st5[31]), .b(st5[45]), .y(st6[45]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa46 (.a(st5[31]), .b(st5[46]), .y(st6[46]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa47 (.a(st5[31]), .b(st5[47]), .y(st6[47]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa48 (.a(st5[31]), .b(st5[48]), .y(st6[48]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa49 (.a(st5[31]), .b(st5[49]), .y(st6[49]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa50 (.a(st5[31]), .b(st5[50]), .y(st6[50]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa51 (.a(st5[31]), .b(st5[51]), .y(st6[51]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa52 (.a(st5[31]), .b(st5[52]), .y(st6[52]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa53 (.a(st5[31]), .b(st5[53]), .y(st6[53]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa54 (.a(st5[31]), .b(st5[54]), .y(st6[54]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa55 (.a(st5[31]), .b(st5[55]), .y(st6[55]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa56 (.a(st5[31]), .b(st5[56]), .y(st6[56]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa57 (.a(st5[31]), .b(st5[57]), .y(st6[57]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa58 (.a(st5[31]), .b(st5[58]), .y(st6[58]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa59 (.a(st5[31]), .b(st5[59]), .y(st6[59]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa60 (.a(st5[31]), .b(st5[60]), .y(st6[60]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa61 (.a(st5[31]), .b(st5[61]), .y(st6[61]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa62 (.a(st5[31]), .b(st5[62]), .y(st6[62]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa63 (.a(st5[31]), .b(st5[63]), .y(st6[63]));
assign st6[64]  = {1'b0, st5[64]};
assign st6[65]  = {1'b0, st5[65]};
assign st6[66]  = {1'b0, st5[66]};
assign st6[67]  = {1'b0, st5[67]};
assign st6[68]  = {1'b0, st5[68]};
assign st6[69]  = {1'b0, st5[69]};
assign st6[70]  = {1'b0, st5[70]};
assign st6[71]  = {1'b0, st5[71]};
assign st6[72]  = {1'b0, st5[72]};
assign st6[73]  = {1'b0, st5[73]};
assign st6[74]  = {1'b0, st5[74]};
assign st6[75]  = {1'b0, st5[75]};
assign st6[76]  = {1'b0, st5[76]};
assign st6[77]  = {1'b0, st5[77]};
assign st6[78]  = {1'b0, st5[78]};
assign st6[79]  = {1'b0, st5[79]};
assign st6[80]  = {1'b0, st5[80]};
assign st6[81]  = {1'b0, st5[81]};
assign st6[82]  = {1'b0, st5[82]};
assign st6[83]  = {1'b0, st5[83]};
assign st6[84]  = {1'b0, st5[84]};
assign st6[85]  = {1'b0, st5[85]};
assign st6[86]  = {1'b0, st5[86]};
assign st6[87]  = {1'b0, st5[87]};
assign st6[88]  = {1'b0, st5[88]};
assign st6[89]  = {1'b0, st5[89]};
assign st6[90]  = {1'b0, st5[90]};
assign st6[91]  = {1'b0, st5[91]};
assign st6[92]  = {1'b0, st5[92]};
assign st6[93]  = {1'b0, st5[93]};
assign st6[94]  = {1'b0, st5[94]};
assign st6[95]  = {1'b0, st5[95]};
NodeAdder #(.WORD_WIDTH(6)) st6_pa96 (.a(st5[95]), .b(st5[96]), .y(st6[96]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa97 (.a(st5[95]), .b(st5[97]), .y(st6[97]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa98 (.a(st5[95]), .b(st5[98]), .y(st6[98]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa99 (.a(st5[95]), .b(st5[99]), .y(st6[99]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa100 (.a(st5[95]), .b(st5[100]), .y(st6[100]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa101 (.a(st5[95]), .b(st5[101]), .y(st6[101]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa102 (.a(st5[95]), .b(st5[102]), .y(st6[102]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa103 (.a(st5[95]), .b(st5[103]), .y(st6[103]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa104 (.a(st5[95]), .b(st5[104]), .y(st6[104]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa105 (.a(st5[95]), .b(st5[105]), .y(st6[105]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa106 (.a(st5[95]), .b(st5[106]), .y(st6[106]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa107 (.a(st5[95]), .b(st5[107]), .y(st6[107]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa108 (.a(st5[95]), .b(st5[108]), .y(st6[108]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa109 (.a(st5[95]), .b(st5[109]), .y(st6[109]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa110 (.a(st5[95]), .b(st5[110]), .y(st6[110]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa111 (.a(st5[95]), .b(st5[111]), .y(st6[111]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa112 (.a(st5[95]), .b(st5[112]), .y(st6[112]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa113 (.a(st5[95]), .b(st5[113]), .y(st6[113]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa114 (.a(st5[95]), .b(st5[114]), .y(st6[114]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa115 (.a(st5[95]), .b(st5[115]), .y(st6[115]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa116 (.a(st5[95]), .b(st5[116]), .y(st6[116]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa117 (.a(st5[95]), .b(st5[117]), .y(st6[117]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa118 (.a(st5[95]), .b(st5[118]), .y(st6[118]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa119 (.a(st5[95]), .b(st5[119]), .y(st6[119]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa120 (.a(st5[95]), .b(st5[120]), .y(st6[120]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa121 (.a(st5[95]), .b(st5[121]), .y(st6[121]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa122 (.a(st5[95]), .b(st5[122]), .y(st6[122]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa123 (.a(st5[95]), .b(st5[123]), .y(st6[123]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa124 (.a(st5[95]), .b(st5[124]), .y(st6[124]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa125 (.a(st5[95]), .b(st5[125]), .y(st6[125]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa126 (.a(st5[95]), .b(st5[126]), .y(st6[126]));
NodeAdder #(.WORD_WIDTH(6)) st6_pa127 (.a(st5[95]), .b(st5[127]), .y(st6[127]));



// Stage 7
wire [7:0] st7 [0:127];

assign st7[0]  = {1'b0, st6[0]};
assign st7[1]  = {1'b0, st6[1]};
assign st7[2]  = {1'b0, st6[2]};
assign st7[3]  = {1'b0, st6[3]};
assign st7[4]  = {1'b0, st6[4]};
assign st7[5]  = {1'b0, st6[5]};
assign st7[6]  = {1'b0, st6[6]};
assign st7[7]  = {1'b0, st6[7]};
assign st7[8]  = {1'b0, st6[8]};
assign st7[9]  = {1'b0, st6[9]};
assign st7[10]  = {1'b0, st6[10]};
assign st7[11]  = {1'b0, st6[11]};
assign st7[12]  = {1'b0, st6[12]};
assign st7[13]  = {1'b0, st6[13]};
assign st7[14]  = {1'b0, st6[14]};
assign st7[15]  = {1'b0, st6[15]};
assign st7[16]  = {1'b0, st6[16]};
assign st7[17]  = {1'b0, st6[17]};
assign st7[18]  = {1'b0, st6[18]};
assign st7[19]  = {1'b0, st6[19]};
assign st7[20]  = {1'b0, st6[20]};
assign st7[21]  = {1'b0, st6[21]};
assign st7[22]  = {1'b0, st6[22]};
assign st7[23]  = {1'b0, st6[23]};
assign st7[24]  = {1'b0, st6[24]};
assign st7[25]  = {1'b0, st6[25]};
assign st7[26]  = {1'b0, st6[26]};
assign st7[27]  = {1'b0, st6[27]};
assign st7[28]  = {1'b0, st6[28]};
assign st7[29]  = {1'b0, st6[29]};
assign st7[30]  = {1'b0, st6[30]};
assign st7[31]  = {1'b0, st6[31]};
assign st7[32]  = {1'b0, st6[32]};
assign st7[33]  = {1'b0, st6[33]};
assign st7[34]  = {1'b0, st6[34]};
assign st7[35]  = {1'b0, st6[35]};
assign st7[36]  = {1'b0, st6[36]};
assign st7[37]  = {1'b0, st6[37]};
assign st7[38]  = {1'b0, st6[38]};
assign st7[39]  = {1'b0, st6[39]};
assign st7[40]  = {1'b0, st6[40]};
assign st7[41]  = {1'b0, st6[41]};
assign st7[42]  = {1'b0, st6[42]};
assign st7[43]  = {1'b0, st6[43]};
assign st7[44]  = {1'b0, st6[44]};
assign st7[45]  = {1'b0, st6[45]};
assign st7[46]  = {1'b0, st6[46]};
assign st7[47]  = {1'b0, st6[47]};
assign st7[48]  = {1'b0, st6[48]};
assign st7[49]  = {1'b0, st6[49]};
assign st7[50]  = {1'b0, st6[50]};
assign st7[51]  = {1'b0, st6[51]};
assign st7[52]  = {1'b0, st6[52]};
assign st7[53]  = {1'b0, st6[53]};
assign st7[54]  = {1'b0, st6[54]};
assign st7[55]  = {1'b0, st6[55]};
assign st7[56]  = {1'b0, st6[56]};
assign st7[57]  = {1'b0, st6[57]};
assign st7[58]  = {1'b0, st6[58]};
assign st7[59]  = {1'b0, st6[59]};
assign st7[60]  = {1'b0, st6[60]};
assign st7[61]  = {1'b0, st6[61]};
assign st7[62]  = {1'b0, st6[62]};
assign st7[63]  = {1'b0, st6[63]};
NodeAdder #(.WORD_WIDTH(7)) st7_pa64 (.a(st6[63]), .b(st6[64]), .y(st7[64]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa65 (.a(st6[63]), .b(st6[65]), .y(st7[65]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa66 (.a(st6[63]), .b(st6[66]), .y(st7[66]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa67 (.a(st6[63]), .b(st6[67]), .y(st7[67]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa68 (.a(st6[63]), .b(st6[68]), .y(st7[68]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa69 (.a(st6[63]), .b(st6[69]), .y(st7[69]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa70 (.a(st6[63]), .b(st6[70]), .y(st7[70]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa71 (.a(st6[63]), .b(st6[71]), .y(st7[71]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa72 (.a(st6[63]), .b(st6[72]), .y(st7[72]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa73 (.a(st6[63]), .b(st6[73]), .y(st7[73]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa74 (.a(st6[63]), .b(st6[74]), .y(st7[74]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa75 (.a(st6[63]), .b(st6[75]), .y(st7[75]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa76 (.a(st6[63]), .b(st6[76]), .y(st7[76]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa77 (.a(st6[63]), .b(st6[77]), .y(st7[77]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa78 (.a(st6[63]), .b(st6[78]), .y(st7[78]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa79 (.a(st6[63]), .b(st6[79]), .y(st7[79]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa80 (.a(st6[63]), .b(st6[80]), .y(st7[80]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa81 (.a(st6[63]), .b(st6[81]), .y(st7[81]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa82 (.a(st6[63]), .b(st6[82]), .y(st7[82]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa83 (.a(st6[63]), .b(st6[83]), .y(st7[83]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa84 (.a(st6[63]), .b(st6[84]), .y(st7[84]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa85 (.a(st6[63]), .b(st6[85]), .y(st7[85]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa86 (.a(st6[63]), .b(st6[86]), .y(st7[86]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa87 (.a(st6[63]), .b(st6[87]), .y(st7[87]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa88 (.a(st6[63]), .b(st6[88]), .y(st7[88]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa89 (.a(st6[63]), .b(st6[89]), .y(st7[89]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa90 (.a(st6[63]), .b(st6[90]), .y(st7[90]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa91 (.a(st6[63]), .b(st6[91]), .y(st7[91]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa92 (.a(st6[63]), .b(st6[92]), .y(st7[92]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa93 (.a(st6[63]), .b(st6[93]), .y(st7[93]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa94 (.a(st6[63]), .b(st6[94]), .y(st7[94]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa95 (.a(st6[63]), .b(st6[95]), .y(st7[95]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa96 (.a(st6[63]), .b(st6[96]), .y(st7[96]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa97 (.a(st6[63]), .b(st6[97]), .y(st7[97]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa98 (.a(st6[63]), .b(st6[98]), .y(st7[98]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa99 (.a(st6[63]), .b(st6[99]), .y(st7[99]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa100 (.a(st6[63]), .b(st6[100]), .y(st7[100]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa101 (.a(st6[63]), .b(st6[101]), .y(st7[101]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa102 (.a(st6[63]), .b(st6[102]), .y(st7[102]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa103 (.a(st6[63]), .b(st6[103]), .y(st7[103]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa104 (.a(st6[63]), .b(st6[104]), .y(st7[104]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa105 (.a(st6[63]), .b(st6[105]), .y(st7[105]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa106 (.a(st6[63]), .b(st6[106]), .y(st7[106]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa107 (.a(st6[63]), .b(st6[107]), .y(st7[107]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa108 (.a(st6[63]), .b(st6[108]), .y(st7[108]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa109 (.a(st6[63]), .b(st6[109]), .y(st7[109]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa110 (.a(st6[63]), .b(st6[110]), .y(st7[110]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa111 (.a(st6[63]), .b(st6[111]), .y(st7[111]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa112 (.a(st6[63]), .b(st6[112]), .y(st7[112]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa113 (.a(st6[63]), .b(st6[113]), .y(st7[113]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa114 (.a(st6[63]), .b(st6[114]), .y(st7[114]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa115 (.a(st6[63]), .b(st6[115]), .y(st7[115]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa116 (.a(st6[63]), .b(st6[116]), .y(st7[116]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa117 (.a(st6[63]), .b(st6[117]), .y(st7[117]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa118 (.a(st6[63]), .b(st6[118]), .y(st7[118]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa119 (.a(st6[63]), .b(st6[119]), .y(st7[119]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa120 (.a(st6[63]), .b(st6[120]), .y(st7[120]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa121 (.a(st6[63]), .b(st6[121]), .y(st7[121]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa122 (.a(st6[63]), .b(st6[122]), .y(st7[122]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa123 (.a(st6[63]), .b(st6[123]), .y(st7[123]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa124 (.a(st6[63]), .b(st6[124]), .y(st7[124]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa125 (.a(st6[63]), .b(st6[125]), .y(st7[125]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa126 (.a(st6[63]), .b(st6[126]), .y(st7[126]));
NodeAdder #(.WORD_WIDTH(7)) st7_pa127 (.a(st6[63]), .b(st6[127]), .y(st7[127]));


// Output link
assign psum[7:0] = st7[0];
assign psum[15:8] = st7[1];
assign psum[23:16] = st7[2];
assign psum[31:24] = st7[3];
assign psum[39:32] = st7[4];
assign psum[47:40] = st7[5];
assign psum[55:48] = st7[6];
assign psum[63:56] = st7[7];
assign psum[71:64] = st7[8];
assign psum[79:72] = st7[9];
assign psum[87:80] = st7[10];
assign psum[95:88] = st7[11];
assign psum[103:96] = st7[12];
assign psum[111:104] = st7[13];
assign psum[119:112] = st7[14];
assign psum[127:120] = st7[15];
assign psum[135:128] = st7[16];
assign psum[143:136] = st7[17];
assign psum[151:144] = st7[18];
assign psum[159:152] = st7[19];
assign psum[167:160] = st7[20];
assign psum[175:168] = st7[21];
assign psum[183:176] = st7[22];
assign psum[191:184] = st7[23];
assign psum[199:192] = st7[24];
assign psum[207:200] = st7[25];
assign psum[215:208] = st7[26];
assign psum[223:216] = st7[27];
assign psum[231:224] = st7[28];
assign psum[239:232] = st7[29];
assign psum[247:240] = st7[30];
assign psum[255:248] = st7[31];
assign psum[263:256] = st7[32];
assign psum[271:264] = st7[33];
assign psum[279:272] = st7[34];
assign psum[287:280] = st7[35];
assign psum[295:288] = st7[36];
assign psum[303:296] = st7[37];
assign psum[311:304] = st7[38];
assign psum[319:312] = st7[39];
assign psum[327:320] = st7[40];
assign psum[335:328] = st7[41];
assign psum[343:336] = st7[42];
assign psum[351:344] = st7[43];
assign psum[359:352] = st7[44];
assign psum[367:360] = st7[45];
assign psum[375:368] = st7[46];
assign psum[383:376] = st7[47];
assign psum[391:384] = st7[48];
assign psum[399:392] = st7[49];
assign psum[407:400] = st7[50];
assign psum[415:408] = st7[51];
assign psum[423:416] = st7[52];
assign psum[431:424] = st7[53];
assign psum[439:432] = st7[54];
assign psum[447:440] = st7[55];
assign psum[455:448] = st7[56];
assign psum[463:456] = st7[57];
assign psum[471:464] = st7[58];
assign psum[479:472] = st7[59];
assign psum[487:480] = st7[60];
assign psum[495:488] = st7[61];
assign psum[503:496] = st7[62];
assign psum[511:504] = st7[63];
assign psum[519:512] = st7[64];
assign psum[527:520] = st7[65];
assign psum[535:528] = st7[66];
assign psum[543:536] = st7[67];
assign psum[551:544] = st7[68];
assign psum[559:552] = st7[69];
assign psum[567:560] = st7[70];
assign psum[575:568] = st7[71];
assign psum[583:576] = st7[72];
assign psum[591:584] = st7[73];
assign psum[599:592] = st7[74];
assign psum[607:600] = st7[75];
assign psum[615:608] = st7[76];
assign psum[623:616] = st7[77];
assign psum[631:624] = st7[78];
assign psum[639:632] = st7[79];
assign psum[647:640] = st7[80];
assign psum[655:648] = st7[81];
assign psum[663:656] = st7[82];
assign psum[671:664] = st7[83];
assign psum[679:672] = st7[84];
assign psum[687:680] = st7[85];
assign psum[695:688] = st7[86];
assign psum[703:696] = st7[87];
assign psum[711:704] = st7[88];
assign psum[719:712] = st7[89];
assign psum[727:720] = st7[90];
assign psum[735:728] = st7[91];
assign psum[743:736] = st7[92];
assign psum[751:744] = st7[93];
assign psum[759:752] = st7[94];
assign psum[767:760] = st7[95];
assign psum[775:768] = st7[96];
assign psum[783:776] = st7[97];
assign psum[791:784] = st7[98];
assign psum[799:792] = st7[99];
assign psum[807:800] = st7[100];
assign psum[815:808] = st7[101];
assign psum[823:816] = st7[102];
assign psum[831:824] = st7[103];
assign psum[839:832] = st7[104];
assign psum[847:840] = st7[105];
assign psum[855:848] = st7[106];
assign psum[863:856] = st7[107];
assign psum[871:864] = st7[108];
assign psum[879:872] = st7[109];
assign psum[887:880] = st7[110];
assign psum[895:888] = st7[111];
assign psum[903:896] = st7[112];
assign psum[911:904] = st7[113];
assign psum[919:912] = st7[114];
assign psum[927:920] = st7[115];
assign psum[935:928] = st7[116];
assign psum[943:936] = st7[117];
assign psum[951:944] = st7[118];
assign psum[959:952] = st7[119];
assign psum[967:960] = st7[120];
assign psum[975:968] = st7[121];
assign psum[983:976] = st7[122];
assign psum[991:984] = st7[123];
assign psum[999:992] = st7[124];
assign psum[1007:1000] = st7[125];
assign psum[1015:1008] = st7[126];
assign psum[1023:1016] = st7[127];

endmodule