module RedundancyController (
    input clk,
    output out,
);
    
endmodule