module BCShifter128 #(  // Bubble-Collapsing Shifter
    parameter WORD_WIDTH    = 8,
    parameter DIST_WIDTH    = 7,
    parameter MAX_LIFM_RSIZ = 3
) (
    input [1023:0] psum,
    input [127:0]  mask,

    input [128*WORD_WIDTH-1:0]               lifm_line,
    input [128*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] mt_line,

    output [128*WORD_WIDTH-1:0]               lifm_comp,
    output [128*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] mt_comp
);

genvar line_idx;  // line index iterator

// Generate array connected with input and output ports
wire [WORD_WIDTH-1:0]               lifm_line_arr [0:127];
wire [DIST_WIDTH*MAX_LIFM_RSIZ-1:0] mt_line_arr   [0:127];

reg [WORD_WIDTH-1:0]               lifm_comp_arr [0:127];
reg [DIST_WIDTH*MAX_LIFM_RSIZ-1:0] mt_comp_arr   [0:127];

generate
    for (line_idx = 0; line_idx < 128; line_idx = line_idx+1) begin
        assign lifm_line_arr[line_idx] = lifm_line[WORD_WIDTH*line_idx+:WORD_WIDTH];
        assign mt_line_arr[line_idx] = mt_line[DIST_WIDTH*MAX_LIFM_RSIZ*line_idx+:DIST_WIDTH*MAX_LIFM_RSIZ];
        assign lifm_comp[WORD_WIDTH*line_idx+:WORD_WIDTH] = lifm_comp_arr[line_idx];
        assign mt_comp[DIST_WIDTH*MAX_LIFM_RSIZ*line_idx+:IST_WIDTH*MAX_LIFM_RSIZ] = mt_comp_arr[line_idx];
    end
endgenerate


// Shifter 2
wire [2*WORD_WIDTH-1:0] i_lifm_l2;
wire [2*WORD_WIDTH-1:0] o_lifm_l2;
wire [2*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l2;
wire [2*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l2;
wire [1:0] stride_l2;

assign i_lifm_l2 = {lifm_line_arr[1], 1*WORD_WIDTH'b0};
assign i_mt_l2 = {mt_line_arr[1], 1*WORD_WIDTH'b0};
assign stride_l2 = psum_arr[1][1:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(2), .NUMEL_LOG(2)
) vs_lifm_2 (
    .i_vec(i_lifm_l2), .stride(stride_l2), .o_vec(o_lifm_l2)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(2), .NUMEL_LOG(2)
) vs_mt_2 (
    .i_vec(i_mt_l2), .stride(stride_l2), .o_vec(o_mt_l2)
);

// Shifter 3
wire [3*WORD_WIDTH-1:0] i_lifm_l3;
wire [3*WORD_WIDTH-1:0] o_lifm_l3;
wire [3*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l3;
wire [3*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l3;
wire [1:0] stride_l3;

assign i_lifm_l3 = {lifm_line_arr[2], 2*WORD_WIDTH'b0};
assign i_mt_l3 = {mt_line_arr[2], 2*WORD_WIDTH'b0};
assign stride_l3 = psum_arr[2][1:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(3), .NUMEL_LOG(2)
) vs_lifm_3 (
    .i_vec(i_lifm_l3), .stride(stride_l3), .o_vec(o_lifm_l3)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(3), .NUMEL_LOG(2)
) vs_mt_3 (
    .i_vec(i_mt_l3), .stride(stride_l3), .o_vec(o_mt_l3)
);

// Shifter 4
wire [4*WORD_WIDTH-1:0] i_lifm_l4;
wire [4*WORD_WIDTH-1:0] o_lifm_l4;
wire [4*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l4;
wire [4*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l4;
wire [2:0] stride_l4;

assign i_lifm_l4 = {lifm_line_arr[3], 3*WORD_WIDTH'b0};
assign i_mt_l4 = {mt_line_arr[3], 3*WORD_WIDTH'b0};
assign stride_l4 = psum_arr[3][2:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(4), .NUMEL_LOG(3)
) vs_lifm_4 (
    .i_vec(i_lifm_l4), .stride(stride_l4), .o_vec(o_lifm_l4)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(4), .NUMEL_LOG(3)
) vs_mt_4 (
    .i_vec(i_mt_l4), .stride(stride_l4), .o_vec(o_mt_l4)
);

// Shifter 5
wire [5*WORD_WIDTH-1:0] i_lifm_l5;
wire [5*WORD_WIDTH-1:0] o_lifm_l5;
wire [5*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l5;
wire [5*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l5;
wire [2:0] stride_l5;

assign i_lifm_l5 = {lifm_line_arr[4], 4*WORD_WIDTH'b0};
assign i_mt_l5 = {mt_line_arr[4], 4*WORD_WIDTH'b0};
assign stride_l5 = psum_arr[4][2:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(5), .NUMEL_LOG(3)
) vs_lifm_5 (
    .i_vec(i_lifm_l5), .stride(stride_l5), .o_vec(o_lifm_l5)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(5), .NUMEL_LOG(3)
) vs_mt_5 (
    .i_vec(i_mt_l5), .stride(stride_l5), .o_vec(o_mt_l5)
);

// Shifter 6
wire [6*WORD_WIDTH-1:0] i_lifm_l6;
wire [6*WORD_WIDTH-1:0] o_lifm_l6;
wire [6*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l6;
wire [6*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l6;
wire [2:0] stride_l6;

assign i_lifm_l6 = {lifm_line_arr[5], 5*WORD_WIDTH'b0};
assign i_mt_l6 = {mt_line_arr[5], 5*WORD_WIDTH'b0};
assign stride_l6 = psum_arr[5][2:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(6), .NUMEL_LOG(3)
) vs_lifm_6 (
    .i_vec(i_lifm_l6), .stride(stride_l6), .o_vec(o_lifm_l6)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(6), .NUMEL_LOG(3)
) vs_mt_6 (
    .i_vec(i_mt_l6), .stride(stride_l6), .o_vec(o_mt_l6)
);

// Shifter 7
wire [7*WORD_WIDTH-1:0] i_lifm_l7;
wire [7*WORD_WIDTH-1:0] o_lifm_l7;
wire [7*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l7;
wire [7*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l7;
wire [2:0] stride_l7;

assign i_lifm_l7 = {lifm_line_arr[6], 6*WORD_WIDTH'b0};
assign i_mt_l7 = {mt_line_arr[6], 6*WORD_WIDTH'b0};
assign stride_l7 = psum_arr[6][2:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(7), .NUMEL_LOG(3)
) vs_lifm_7 (
    .i_vec(i_lifm_l7), .stride(stride_l7), .o_vec(o_lifm_l7)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(7), .NUMEL_LOG(3)
) vs_mt_7 (
    .i_vec(i_mt_l7), .stride(stride_l7), .o_vec(o_mt_l7)
);

// Shifter 8
wire [8*WORD_WIDTH-1:0] i_lifm_l8;
wire [8*WORD_WIDTH-1:0] o_lifm_l8;
wire [8*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l8;
wire [8*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l8;
wire [3:0] stride_l8;

assign i_lifm_l8 = {lifm_line_arr[7], 7*WORD_WIDTH'b0};
assign i_mt_l8 = {mt_line_arr[7], 7*WORD_WIDTH'b0};
assign stride_l8 = psum_arr[7][3:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(8), .NUMEL_LOG(4)
) vs_lifm_8 (
    .i_vec(i_lifm_l8), .stride(stride_l8), .o_vec(o_lifm_l8)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(8), .NUMEL_LOG(4)
) vs_mt_8 (
    .i_vec(i_mt_l8), .stride(stride_l8), .o_vec(o_mt_l8)
);

// Shifter 9
wire [9*WORD_WIDTH-1:0] i_lifm_l9;
wire [9*WORD_WIDTH-1:0] o_lifm_l9;
wire [9*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l9;
wire [9*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l9;
wire [3:0] stride_l9;

assign i_lifm_l9 = {lifm_line_arr[8], 8*WORD_WIDTH'b0};
assign i_mt_l9 = {mt_line_arr[8], 8*WORD_WIDTH'b0};
assign stride_l9 = psum_arr[8][3:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(9), .NUMEL_LOG(4)
) vs_lifm_9 (
    .i_vec(i_lifm_l9), .stride(stride_l9), .o_vec(o_lifm_l9)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(9), .NUMEL_LOG(4)
) vs_mt_9 (
    .i_vec(i_mt_l9), .stride(stride_l9), .o_vec(o_mt_l9)
);

// Shifter 10
wire [10*WORD_WIDTH-1:0] i_lifm_l10;
wire [10*WORD_WIDTH-1:0] o_lifm_l10;
wire [10*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l10;
wire [10*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l10;
wire [3:0] stride_l10;

assign i_lifm_l10 = {lifm_line_arr[9], 9*WORD_WIDTH'b0};
assign i_mt_l10 = {mt_line_arr[9], 9*WORD_WIDTH'b0};
assign stride_l10 = psum_arr[9][3:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(10), .NUMEL_LOG(4)
) vs_lifm_10 (
    .i_vec(i_lifm_l10), .stride(stride_l10), .o_vec(o_lifm_l10)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(10), .NUMEL_LOG(4)
) vs_mt_10 (
    .i_vec(i_mt_l10), .stride(stride_l10), .o_vec(o_mt_l10)
);

// Shifter 11
wire [11*WORD_WIDTH-1:0] i_lifm_l11;
wire [11*WORD_WIDTH-1:0] o_lifm_l11;
wire [11*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l11;
wire [11*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l11;
wire [3:0] stride_l11;

assign i_lifm_l11 = {lifm_line_arr[10], 10*WORD_WIDTH'b0};
assign i_mt_l11 = {mt_line_arr[10], 10*WORD_WIDTH'b0};
assign stride_l11 = psum_arr[10][3:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(11), .NUMEL_LOG(4)
) vs_lifm_11 (
    .i_vec(i_lifm_l11), .stride(stride_l11), .o_vec(o_lifm_l11)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(11), .NUMEL_LOG(4)
) vs_mt_11 (
    .i_vec(i_mt_l11), .stride(stride_l11), .o_vec(o_mt_l11)
);

// Shifter 12
wire [12*WORD_WIDTH-1:0] i_lifm_l12;
wire [12*WORD_WIDTH-1:0] o_lifm_l12;
wire [12*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l12;
wire [12*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l12;
wire [3:0] stride_l12;

assign i_lifm_l12 = {lifm_line_arr[11], 11*WORD_WIDTH'b0};
assign i_mt_l12 = {mt_line_arr[11], 11*WORD_WIDTH'b0};
assign stride_l12 = psum_arr[11][3:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(12), .NUMEL_LOG(4)
) vs_lifm_12 (
    .i_vec(i_lifm_l12), .stride(stride_l12), .o_vec(o_lifm_l12)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(12), .NUMEL_LOG(4)
) vs_mt_12 (
    .i_vec(i_mt_l12), .stride(stride_l12), .o_vec(o_mt_l12)
);

// Shifter 13
wire [13*WORD_WIDTH-1:0] i_lifm_l13;
wire [13*WORD_WIDTH-1:0] o_lifm_l13;
wire [13*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l13;
wire [13*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l13;
wire [3:0] stride_l13;

assign i_lifm_l13 = {lifm_line_arr[12], 12*WORD_WIDTH'b0};
assign i_mt_l13 = {mt_line_arr[12], 12*WORD_WIDTH'b0};
assign stride_l13 = psum_arr[12][3:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(13), .NUMEL_LOG(4)
) vs_lifm_13 (
    .i_vec(i_lifm_l13), .stride(stride_l13), .o_vec(o_lifm_l13)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(13), .NUMEL_LOG(4)
) vs_mt_13 (
    .i_vec(i_mt_l13), .stride(stride_l13), .o_vec(o_mt_l13)
);

// Shifter 14
wire [14*WORD_WIDTH-1:0] i_lifm_l14;
wire [14*WORD_WIDTH-1:0] o_lifm_l14;
wire [14*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l14;
wire [14*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l14;
wire [3:0] stride_l14;

assign i_lifm_l14 = {lifm_line_arr[13], 13*WORD_WIDTH'b0};
assign i_mt_l14 = {mt_line_arr[13], 13*WORD_WIDTH'b0};
assign stride_l14 = psum_arr[13][3:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(14), .NUMEL_LOG(4)
) vs_lifm_14 (
    .i_vec(i_lifm_l14), .stride(stride_l14), .o_vec(o_lifm_l14)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(14), .NUMEL_LOG(4)
) vs_mt_14 (
    .i_vec(i_mt_l14), .stride(stride_l14), .o_vec(o_mt_l14)
);

// Shifter 15
wire [15*WORD_WIDTH-1:0] i_lifm_l15;
wire [15*WORD_WIDTH-1:0] o_lifm_l15;
wire [15*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l15;
wire [15*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l15;
wire [3:0] stride_l15;

assign i_lifm_l15 = {lifm_line_arr[14], 14*WORD_WIDTH'b0};
assign i_mt_l15 = {mt_line_arr[14], 14*WORD_WIDTH'b0};
assign stride_l15 = psum_arr[14][3:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(15), .NUMEL_LOG(4)
) vs_lifm_15 (
    .i_vec(i_lifm_l15), .stride(stride_l15), .o_vec(o_lifm_l15)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(15), .NUMEL_LOG(4)
) vs_mt_15 (
    .i_vec(i_mt_l15), .stride(stride_l15), .o_vec(o_mt_l15)
);

// Shifter 16
wire [16*WORD_WIDTH-1:0] i_lifm_l16;
wire [16*WORD_WIDTH-1:0] o_lifm_l16;
wire [16*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l16;
wire [16*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l16;
wire [4:0] stride_l16;

assign i_lifm_l16 = {lifm_line_arr[15], 15*WORD_WIDTH'b0};
assign i_mt_l16 = {mt_line_arr[15], 15*WORD_WIDTH'b0};
assign stride_l16 = psum_arr[15][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(16), .NUMEL_LOG(5)
) vs_lifm_16 (
    .i_vec(i_lifm_l16), .stride(stride_l16), .o_vec(o_lifm_l16)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(16), .NUMEL_LOG(5)
) vs_mt_16 (
    .i_vec(i_mt_l16), .stride(stride_l16), .o_vec(o_mt_l16)
);

// Shifter 17
wire [17*WORD_WIDTH-1:0] i_lifm_l17;
wire [17*WORD_WIDTH-1:0] o_lifm_l17;
wire [17*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l17;
wire [17*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l17;
wire [4:0] stride_l17;

assign i_lifm_l17 = {lifm_line_arr[16], 16*WORD_WIDTH'b0};
assign i_mt_l17 = {mt_line_arr[16], 16*WORD_WIDTH'b0};
assign stride_l17 = psum_arr[16][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(17), .NUMEL_LOG(5)
) vs_lifm_17 (
    .i_vec(i_lifm_l17), .stride(stride_l17), .o_vec(o_lifm_l17)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(17), .NUMEL_LOG(5)
) vs_mt_17 (
    .i_vec(i_mt_l17), .stride(stride_l17), .o_vec(o_mt_l17)
);

// Shifter 18
wire [18*WORD_WIDTH-1:0] i_lifm_l18;
wire [18*WORD_WIDTH-1:0] o_lifm_l18;
wire [18*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l18;
wire [18*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l18;
wire [4:0] stride_l18;

assign i_lifm_l18 = {lifm_line_arr[17], 17*WORD_WIDTH'b0};
assign i_mt_l18 = {mt_line_arr[17], 17*WORD_WIDTH'b0};
assign stride_l18 = psum_arr[17][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(18), .NUMEL_LOG(5)
) vs_lifm_18 (
    .i_vec(i_lifm_l18), .stride(stride_l18), .o_vec(o_lifm_l18)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(18), .NUMEL_LOG(5)
) vs_mt_18 (
    .i_vec(i_mt_l18), .stride(stride_l18), .o_vec(o_mt_l18)
);

// Shifter 19
wire [19*WORD_WIDTH-1:0] i_lifm_l19;
wire [19*WORD_WIDTH-1:0] o_lifm_l19;
wire [19*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l19;
wire [19*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l19;
wire [4:0] stride_l19;

assign i_lifm_l19 = {lifm_line_arr[18], 18*WORD_WIDTH'b0};
assign i_mt_l19 = {mt_line_arr[18], 18*WORD_WIDTH'b0};
assign stride_l19 = psum_arr[18][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(19), .NUMEL_LOG(5)
) vs_lifm_19 (
    .i_vec(i_lifm_l19), .stride(stride_l19), .o_vec(o_lifm_l19)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(19), .NUMEL_LOG(5)
) vs_mt_19 (
    .i_vec(i_mt_l19), .stride(stride_l19), .o_vec(o_mt_l19)
);

// Shifter 20
wire [20*WORD_WIDTH-1:0] i_lifm_l20;
wire [20*WORD_WIDTH-1:0] o_lifm_l20;
wire [20*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l20;
wire [20*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l20;
wire [4:0] stride_l20;

assign i_lifm_l20 = {lifm_line_arr[19], 19*WORD_WIDTH'b0};
assign i_mt_l20 = {mt_line_arr[19], 19*WORD_WIDTH'b0};
assign stride_l20 = psum_arr[19][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(20), .NUMEL_LOG(5)
) vs_lifm_20 (
    .i_vec(i_lifm_l20), .stride(stride_l20), .o_vec(o_lifm_l20)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(20), .NUMEL_LOG(5)
) vs_mt_20 (
    .i_vec(i_mt_l20), .stride(stride_l20), .o_vec(o_mt_l20)
);

// Shifter 21
wire [21*WORD_WIDTH-1:0] i_lifm_l21;
wire [21*WORD_WIDTH-1:0] o_lifm_l21;
wire [21*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l21;
wire [21*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l21;
wire [4:0] stride_l21;

assign i_lifm_l21 = {lifm_line_arr[20], 20*WORD_WIDTH'b0};
assign i_mt_l21 = {mt_line_arr[20], 20*WORD_WIDTH'b0};
assign stride_l21 = psum_arr[20][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(21), .NUMEL_LOG(5)
) vs_lifm_21 (
    .i_vec(i_lifm_l21), .stride(stride_l21), .o_vec(o_lifm_l21)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(21), .NUMEL_LOG(5)
) vs_mt_21 (
    .i_vec(i_mt_l21), .stride(stride_l21), .o_vec(o_mt_l21)
);

// Shifter 22
wire [22*WORD_WIDTH-1:0] i_lifm_l22;
wire [22*WORD_WIDTH-1:0] o_lifm_l22;
wire [22*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l22;
wire [22*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l22;
wire [4:0] stride_l22;

assign i_lifm_l22 = {lifm_line_arr[21], 21*WORD_WIDTH'b0};
assign i_mt_l22 = {mt_line_arr[21], 21*WORD_WIDTH'b0};
assign stride_l22 = psum_arr[21][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(22), .NUMEL_LOG(5)
) vs_lifm_22 (
    .i_vec(i_lifm_l22), .stride(stride_l22), .o_vec(o_lifm_l22)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(22), .NUMEL_LOG(5)
) vs_mt_22 (
    .i_vec(i_mt_l22), .stride(stride_l22), .o_vec(o_mt_l22)
);

// Shifter 23
wire [23*WORD_WIDTH-1:0] i_lifm_l23;
wire [23*WORD_WIDTH-1:0] o_lifm_l23;
wire [23*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l23;
wire [23*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l23;
wire [4:0] stride_l23;

assign i_lifm_l23 = {lifm_line_arr[22], 22*WORD_WIDTH'b0};
assign i_mt_l23 = {mt_line_arr[22], 22*WORD_WIDTH'b0};
assign stride_l23 = psum_arr[22][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(23), .NUMEL_LOG(5)
) vs_lifm_23 (
    .i_vec(i_lifm_l23), .stride(stride_l23), .o_vec(o_lifm_l23)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(23), .NUMEL_LOG(5)
) vs_mt_23 (
    .i_vec(i_mt_l23), .stride(stride_l23), .o_vec(o_mt_l23)
);

// Shifter 24
wire [24*WORD_WIDTH-1:0] i_lifm_l24;
wire [24*WORD_WIDTH-1:0] o_lifm_l24;
wire [24*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l24;
wire [24*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l24;
wire [4:0] stride_l24;

assign i_lifm_l24 = {lifm_line_arr[23], 23*WORD_WIDTH'b0};
assign i_mt_l24 = {mt_line_arr[23], 23*WORD_WIDTH'b0};
assign stride_l24 = psum_arr[23][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(24), .NUMEL_LOG(5)
) vs_lifm_24 (
    .i_vec(i_lifm_l24), .stride(stride_l24), .o_vec(o_lifm_l24)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(24), .NUMEL_LOG(5)
) vs_mt_24 (
    .i_vec(i_mt_l24), .stride(stride_l24), .o_vec(o_mt_l24)
);

// Shifter 25
wire [25*WORD_WIDTH-1:0] i_lifm_l25;
wire [25*WORD_WIDTH-1:0] o_lifm_l25;
wire [25*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l25;
wire [25*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l25;
wire [4:0] stride_l25;

assign i_lifm_l25 = {lifm_line_arr[24], 24*WORD_WIDTH'b0};
assign i_mt_l25 = {mt_line_arr[24], 24*WORD_WIDTH'b0};
assign stride_l25 = psum_arr[24][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(25), .NUMEL_LOG(5)
) vs_lifm_25 (
    .i_vec(i_lifm_l25), .stride(stride_l25), .o_vec(o_lifm_l25)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(25), .NUMEL_LOG(5)
) vs_mt_25 (
    .i_vec(i_mt_l25), .stride(stride_l25), .o_vec(o_mt_l25)
);

// Shifter 26
wire [26*WORD_WIDTH-1:0] i_lifm_l26;
wire [26*WORD_WIDTH-1:0] o_lifm_l26;
wire [26*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l26;
wire [26*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l26;
wire [4:0] stride_l26;

assign i_lifm_l26 = {lifm_line_arr[25], 25*WORD_WIDTH'b0};
assign i_mt_l26 = {mt_line_arr[25], 25*WORD_WIDTH'b0};
assign stride_l26 = psum_arr[25][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(26), .NUMEL_LOG(5)
) vs_lifm_26 (
    .i_vec(i_lifm_l26), .stride(stride_l26), .o_vec(o_lifm_l26)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(26), .NUMEL_LOG(5)
) vs_mt_26 (
    .i_vec(i_mt_l26), .stride(stride_l26), .o_vec(o_mt_l26)
);

// Shifter 27
wire [27*WORD_WIDTH-1:0] i_lifm_l27;
wire [27*WORD_WIDTH-1:0] o_lifm_l27;
wire [27*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l27;
wire [27*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l27;
wire [4:0] stride_l27;

assign i_lifm_l27 = {lifm_line_arr[26], 26*WORD_WIDTH'b0};
assign i_mt_l27 = {mt_line_arr[26], 26*WORD_WIDTH'b0};
assign stride_l27 = psum_arr[26][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(27), .NUMEL_LOG(5)
) vs_lifm_27 (
    .i_vec(i_lifm_l27), .stride(stride_l27), .o_vec(o_lifm_l27)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(27), .NUMEL_LOG(5)
) vs_mt_27 (
    .i_vec(i_mt_l27), .stride(stride_l27), .o_vec(o_mt_l27)
);

// Shifter 28
wire [28*WORD_WIDTH-1:0] i_lifm_l28;
wire [28*WORD_WIDTH-1:0] o_lifm_l28;
wire [28*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l28;
wire [28*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l28;
wire [4:0] stride_l28;

assign i_lifm_l28 = {lifm_line_arr[27], 27*WORD_WIDTH'b0};
assign i_mt_l28 = {mt_line_arr[27], 27*WORD_WIDTH'b0};
assign stride_l28 = psum_arr[27][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(28), .NUMEL_LOG(5)
) vs_lifm_28 (
    .i_vec(i_lifm_l28), .stride(stride_l28), .o_vec(o_lifm_l28)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(28), .NUMEL_LOG(5)
) vs_mt_28 (
    .i_vec(i_mt_l28), .stride(stride_l28), .o_vec(o_mt_l28)
);

// Shifter 29
wire [29*WORD_WIDTH-1:0] i_lifm_l29;
wire [29*WORD_WIDTH-1:0] o_lifm_l29;
wire [29*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l29;
wire [29*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l29;
wire [4:0] stride_l29;

assign i_lifm_l29 = {lifm_line_arr[28], 28*WORD_WIDTH'b0};
assign i_mt_l29 = {mt_line_arr[28], 28*WORD_WIDTH'b0};
assign stride_l29 = psum_arr[28][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(29), .NUMEL_LOG(5)
) vs_lifm_29 (
    .i_vec(i_lifm_l29), .stride(stride_l29), .o_vec(o_lifm_l29)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(29), .NUMEL_LOG(5)
) vs_mt_29 (
    .i_vec(i_mt_l29), .stride(stride_l29), .o_vec(o_mt_l29)
);

// Shifter 30
wire [30*WORD_WIDTH-1:0] i_lifm_l30;
wire [30*WORD_WIDTH-1:0] o_lifm_l30;
wire [30*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l30;
wire [30*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l30;
wire [4:0] stride_l30;

assign i_lifm_l30 = {lifm_line_arr[29], 29*WORD_WIDTH'b0};
assign i_mt_l30 = {mt_line_arr[29], 29*WORD_WIDTH'b0};
assign stride_l30 = psum_arr[29][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(30), .NUMEL_LOG(5)
) vs_lifm_30 (
    .i_vec(i_lifm_l30), .stride(stride_l30), .o_vec(o_lifm_l30)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(30), .NUMEL_LOG(5)
) vs_mt_30 (
    .i_vec(i_mt_l30), .stride(stride_l30), .o_vec(o_mt_l30)
);

// Shifter 31
wire [31*WORD_WIDTH-1:0] i_lifm_l31;
wire [31*WORD_WIDTH-1:0] o_lifm_l31;
wire [31*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l31;
wire [31*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l31;
wire [4:0] stride_l31;

assign i_lifm_l31 = {lifm_line_arr[30], 30*WORD_WIDTH'b0};
assign i_mt_l31 = {mt_line_arr[30], 30*WORD_WIDTH'b0};
assign stride_l31 = psum_arr[30][4:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(31), .NUMEL_LOG(5)
) vs_lifm_31 (
    .i_vec(i_lifm_l31), .stride(stride_l31), .o_vec(o_lifm_l31)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(31), .NUMEL_LOG(5)
) vs_mt_31 (
    .i_vec(i_mt_l31), .stride(stride_l31), .o_vec(o_mt_l31)
);

// Shifter 32
wire [32*WORD_WIDTH-1:0] i_lifm_l32;
wire [32*WORD_WIDTH-1:0] o_lifm_l32;
wire [32*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l32;
wire [32*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l32;
wire [5:0] stride_l32;

assign i_lifm_l32 = {lifm_line_arr[31], 31*WORD_WIDTH'b0};
assign i_mt_l32 = {mt_line_arr[31], 31*WORD_WIDTH'b0};
assign stride_l32 = psum_arr[31][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(32), .NUMEL_LOG(6)
) vs_lifm_32 (
    .i_vec(i_lifm_l32), .stride(stride_l32), .o_vec(o_lifm_l32)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(32), .NUMEL_LOG(6)
) vs_mt_32 (
    .i_vec(i_mt_l32), .stride(stride_l32), .o_vec(o_mt_l32)
);

// Shifter 33
wire [33*WORD_WIDTH-1:0] i_lifm_l33;
wire [33*WORD_WIDTH-1:0] o_lifm_l33;
wire [33*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l33;
wire [33*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l33;
wire [5:0] stride_l33;

assign i_lifm_l33 = {lifm_line_arr[32], 32*WORD_WIDTH'b0};
assign i_mt_l33 = {mt_line_arr[32], 32*WORD_WIDTH'b0};
assign stride_l33 = psum_arr[32][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(33), .NUMEL_LOG(6)
) vs_lifm_33 (
    .i_vec(i_lifm_l33), .stride(stride_l33), .o_vec(o_lifm_l33)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(33), .NUMEL_LOG(6)
) vs_mt_33 (
    .i_vec(i_mt_l33), .stride(stride_l33), .o_vec(o_mt_l33)
);

// Shifter 34
wire [34*WORD_WIDTH-1:0] i_lifm_l34;
wire [34*WORD_WIDTH-1:0] o_lifm_l34;
wire [34*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l34;
wire [34*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l34;
wire [5:0] stride_l34;

assign i_lifm_l34 = {lifm_line_arr[33], 33*WORD_WIDTH'b0};
assign i_mt_l34 = {mt_line_arr[33], 33*WORD_WIDTH'b0};
assign stride_l34 = psum_arr[33][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(34), .NUMEL_LOG(6)
) vs_lifm_34 (
    .i_vec(i_lifm_l34), .stride(stride_l34), .o_vec(o_lifm_l34)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(34), .NUMEL_LOG(6)
) vs_mt_34 (
    .i_vec(i_mt_l34), .stride(stride_l34), .o_vec(o_mt_l34)
);

// Shifter 35
wire [35*WORD_WIDTH-1:0] i_lifm_l35;
wire [35*WORD_WIDTH-1:0] o_lifm_l35;
wire [35*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l35;
wire [35*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l35;
wire [5:0] stride_l35;

assign i_lifm_l35 = {lifm_line_arr[34], 34*WORD_WIDTH'b0};
assign i_mt_l35 = {mt_line_arr[34], 34*WORD_WIDTH'b0};
assign stride_l35 = psum_arr[34][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(35), .NUMEL_LOG(6)
) vs_lifm_35 (
    .i_vec(i_lifm_l35), .stride(stride_l35), .o_vec(o_lifm_l35)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(35), .NUMEL_LOG(6)
) vs_mt_35 (
    .i_vec(i_mt_l35), .stride(stride_l35), .o_vec(o_mt_l35)
);

// Shifter 36
wire [36*WORD_WIDTH-1:0] i_lifm_l36;
wire [36*WORD_WIDTH-1:0] o_lifm_l36;
wire [36*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l36;
wire [36*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l36;
wire [5:0] stride_l36;

assign i_lifm_l36 = {lifm_line_arr[35], 35*WORD_WIDTH'b0};
assign i_mt_l36 = {mt_line_arr[35], 35*WORD_WIDTH'b0};
assign stride_l36 = psum_arr[35][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(36), .NUMEL_LOG(6)
) vs_lifm_36 (
    .i_vec(i_lifm_l36), .stride(stride_l36), .o_vec(o_lifm_l36)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(36), .NUMEL_LOG(6)
) vs_mt_36 (
    .i_vec(i_mt_l36), .stride(stride_l36), .o_vec(o_mt_l36)
);

// Shifter 37
wire [37*WORD_WIDTH-1:0] i_lifm_l37;
wire [37*WORD_WIDTH-1:0] o_lifm_l37;
wire [37*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l37;
wire [37*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l37;
wire [5:0] stride_l37;

assign i_lifm_l37 = {lifm_line_arr[36], 36*WORD_WIDTH'b0};
assign i_mt_l37 = {mt_line_arr[36], 36*WORD_WIDTH'b0};
assign stride_l37 = psum_arr[36][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(37), .NUMEL_LOG(6)
) vs_lifm_37 (
    .i_vec(i_lifm_l37), .stride(stride_l37), .o_vec(o_lifm_l37)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(37), .NUMEL_LOG(6)
) vs_mt_37 (
    .i_vec(i_mt_l37), .stride(stride_l37), .o_vec(o_mt_l37)
);

// Shifter 38
wire [38*WORD_WIDTH-1:0] i_lifm_l38;
wire [38*WORD_WIDTH-1:0] o_lifm_l38;
wire [38*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l38;
wire [38*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l38;
wire [5:0] stride_l38;

assign i_lifm_l38 = {lifm_line_arr[37], 37*WORD_WIDTH'b0};
assign i_mt_l38 = {mt_line_arr[37], 37*WORD_WIDTH'b0};
assign stride_l38 = psum_arr[37][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(38), .NUMEL_LOG(6)
) vs_lifm_38 (
    .i_vec(i_lifm_l38), .stride(stride_l38), .o_vec(o_lifm_l38)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(38), .NUMEL_LOG(6)
) vs_mt_38 (
    .i_vec(i_mt_l38), .stride(stride_l38), .o_vec(o_mt_l38)
);

// Shifter 39
wire [39*WORD_WIDTH-1:0] i_lifm_l39;
wire [39*WORD_WIDTH-1:0] o_lifm_l39;
wire [39*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l39;
wire [39*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l39;
wire [5:0] stride_l39;

assign i_lifm_l39 = {lifm_line_arr[38], 38*WORD_WIDTH'b0};
assign i_mt_l39 = {mt_line_arr[38], 38*WORD_WIDTH'b0};
assign stride_l39 = psum_arr[38][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(39), .NUMEL_LOG(6)
) vs_lifm_39 (
    .i_vec(i_lifm_l39), .stride(stride_l39), .o_vec(o_lifm_l39)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(39), .NUMEL_LOG(6)
) vs_mt_39 (
    .i_vec(i_mt_l39), .stride(stride_l39), .o_vec(o_mt_l39)
);

// Shifter 40
wire [40*WORD_WIDTH-1:0] i_lifm_l40;
wire [40*WORD_WIDTH-1:0] o_lifm_l40;
wire [40*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l40;
wire [40*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l40;
wire [5:0] stride_l40;

assign i_lifm_l40 = {lifm_line_arr[39], 39*WORD_WIDTH'b0};
assign i_mt_l40 = {mt_line_arr[39], 39*WORD_WIDTH'b0};
assign stride_l40 = psum_arr[39][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(40), .NUMEL_LOG(6)
) vs_lifm_40 (
    .i_vec(i_lifm_l40), .stride(stride_l40), .o_vec(o_lifm_l40)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(40), .NUMEL_LOG(6)
) vs_mt_40 (
    .i_vec(i_mt_l40), .stride(stride_l40), .o_vec(o_mt_l40)
);

// Shifter 41
wire [41*WORD_WIDTH-1:0] i_lifm_l41;
wire [41*WORD_WIDTH-1:0] o_lifm_l41;
wire [41*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l41;
wire [41*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l41;
wire [5:0] stride_l41;

assign i_lifm_l41 = {lifm_line_arr[40], 40*WORD_WIDTH'b0};
assign i_mt_l41 = {mt_line_arr[40], 40*WORD_WIDTH'b0};
assign stride_l41 = psum_arr[40][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(41), .NUMEL_LOG(6)
) vs_lifm_41 (
    .i_vec(i_lifm_l41), .stride(stride_l41), .o_vec(o_lifm_l41)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(41), .NUMEL_LOG(6)
) vs_mt_41 (
    .i_vec(i_mt_l41), .stride(stride_l41), .o_vec(o_mt_l41)
);

// Shifter 42
wire [42*WORD_WIDTH-1:0] i_lifm_l42;
wire [42*WORD_WIDTH-1:0] o_lifm_l42;
wire [42*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l42;
wire [42*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l42;
wire [5:0] stride_l42;

assign i_lifm_l42 = {lifm_line_arr[41], 41*WORD_WIDTH'b0};
assign i_mt_l42 = {mt_line_arr[41], 41*WORD_WIDTH'b0};
assign stride_l42 = psum_arr[41][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(42), .NUMEL_LOG(6)
) vs_lifm_42 (
    .i_vec(i_lifm_l42), .stride(stride_l42), .o_vec(o_lifm_l42)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(42), .NUMEL_LOG(6)
) vs_mt_42 (
    .i_vec(i_mt_l42), .stride(stride_l42), .o_vec(o_mt_l42)
);

// Shifter 43
wire [43*WORD_WIDTH-1:0] i_lifm_l43;
wire [43*WORD_WIDTH-1:0] o_lifm_l43;
wire [43*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l43;
wire [43*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l43;
wire [5:0] stride_l43;

assign i_lifm_l43 = {lifm_line_arr[42], 42*WORD_WIDTH'b0};
assign i_mt_l43 = {mt_line_arr[42], 42*WORD_WIDTH'b0};
assign stride_l43 = psum_arr[42][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(43), .NUMEL_LOG(6)
) vs_lifm_43 (
    .i_vec(i_lifm_l43), .stride(stride_l43), .o_vec(o_lifm_l43)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(43), .NUMEL_LOG(6)
) vs_mt_43 (
    .i_vec(i_mt_l43), .stride(stride_l43), .o_vec(o_mt_l43)
);

// Shifter 44
wire [44*WORD_WIDTH-1:0] i_lifm_l44;
wire [44*WORD_WIDTH-1:0] o_lifm_l44;
wire [44*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l44;
wire [44*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l44;
wire [5:0] stride_l44;

assign i_lifm_l44 = {lifm_line_arr[43], 43*WORD_WIDTH'b0};
assign i_mt_l44 = {mt_line_arr[43], 43*WORD_WIDTH'b0};
assign stride_l44 = psum_arr[43][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(44), .NUMEL_LOG(6)
) vs_lifm_44 (
    .i_vec(i_lifm_l44), .stride(stride_l44), .o_vec(o_lifm_l44)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(44), .NUMEL_LOG(6)
) vs_mt_44 (
    .i_vec(i_mt_l44), .stride(stride_l44), .o_vec(o_mt_l44)
);

// Shifter 45
wire [45*WORD_WIDTH-1:0] i_lifm_l45;
wire [45*WORD_WIDTH-1:0] o_lifm_l45;
wire [45*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l45;
wire [45*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l45;
wire [5:0] stride_l45;

assign i_lifm_l45 = {lifm_line_arr[44], 44*WORD_WIDTH'b0};
assign i_mt_l45 = {mt_line_arr[44], 44*WORD_WIDTH'b0};
assign stride_l45 = psum_arr[44][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(45), .NUMEL_LOG(6)
) vs_lifm_45 (
    .i_vec(i_lifm_l45), .stride(stride_l45), .o_vec(o_lifm_l45)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(45), .NUMEL_LOG(6)
) vs_mt_45 (
    .i_vec(i_mt_l45), .stride(stride_l45), .o_vec(o_mt_l45)
);

// Shifter 46
wire [46*WORD_WIDTH-1:0] i_lifm_l46;
wire [46*WORD_WIDTH-1:0] o_lifm_l46;
wire [46*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l46;
wire [46*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l46;
wire [5:0] stride_l46;

assign i_lifm_l46 = {lifm_line_arr[45], 45*WORD_WIDTH'b0};
assign i_mt_l46 = {mt_line_arr[45], 45*WORD_WIDTH'b0};
assign stride_l46 = psum_arr[45][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(46), .NUMEL_LOG(6)
) vs_lifm_46 (
    .i_vec(i_lifm_l46), .stride(stride_l46), .o_vec(o_lifm_l46)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(46), .NUMEL_LOG(6)
) vs_mt_46 (
    .i_vec(i_mt_l46), .stride(stride_l46), .o_vec(o_mt_l46)
);

// Shifter 47
wire [47*WORD_WIDTH-1:0] i_lifm_l47;
wire [47*WORD_WIDTH-1:0] o_lifm_l47;
wire [47*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l47;
wire [47*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l47;
wire [5:0] stride_l47;

assign i_lifm_l47 = {lifm_line_arr[46], 46*WORD_WIDTH'b0};
assign i_mt_l47 = {mt_line_arr[46], 46*WORD_WIDTH'b0};
assign stride_l47 = psum_arr[46][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(47), .NUMEL_LOG(6)
) vs_lifm_47 (
    .i_vec(i_lifm_l47), .stride(stride_l47), .o_vec(o_lifm_l47)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(47), .NUMEL_LOG(6)
) vs_mt_47 (
    .i_vec(i_mt_l47), .stride(stride_l47), .o_vec(o_mt_l47)
);

// Shifter 48
wire [48*WORD_WIDTH-1:0] i_lifm_l48;
wire [48*WORD_WIDTH-1:0] o_lifm_l48;
wire [48*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l48;
wire [48*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l48;
wire [5:0] stride_l48;

assign i_lifm_l48 = {lifm_line_arr[47], 47*WORD_WIDTH'b0};
assign i_mt_l48 = {mt_line_arr[47], 47*WORD_WIDTH'b0};
assign stride_l48 = psum_arr[47][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(48), .NUMEL_LOG(6)
) vs_lifm_48 (
    .i_vec(i_lifm_l48), .stride(stride_l48), .o_vec(o_lifm_l48)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(48), .NUMEL_LOG(6)
) vs_mt_48 (
    .i_vec(i_mt_l48), .stride(stride_l48), .o_vec(o_mt_l48)
);

// Shifter 49
wire [49*WORD_WIDTH-1:0] i_lifm_l49;
wire [49*WORD_WIDTH-1:0] o_lifm_l49;
wire [49*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l49;
wire [49*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l49;
wire [5:0] stride_l49;

assign i_lifm_l49 = {lifm_line_arr[48], 48*WORD_WIDTH'b0};
assign i_mt_l49 = {mt_line_arr[48], 48*WORD_WIDTH'b0};
assign stride_l49 = psum_arr[48][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(49), .NUMEL_LOG(6)
) vs_lifm_49 (
    .i_vec(i_lifm_l49), .stride(stride_l49), .o_vec(o_lifm_l49)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(49), .NUMEL_LOG(6)
) vs_mt_49 (
    .i_vec(i_mt_l49), .stride(stride_l49), .o_vec(o_mt_l49)
);

// Shifter 50
wire [50*WORD_WIDTH-1:0] i_lifm_l50;
wire [50*WORD_WIDTH-1:0] o_lifm_l50;
wire [50*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l50;
wire [50*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l50;
wire [5:0] stride_l50;

assign i_lifm_l50 = {lifm_line_arr[49], 49*WORD_WIDTH'b0};
assign i_mt_l50 = {mt_line_arr[49], 49*WORD_WIDTH'b0};
assign stride_l50 = psum_arr[49][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(50), .NUMEL_LOG(6)
) vs_lifm_50 (
    .i_vec(i_lifm_l50), .stride(stride_l50), .o_vec(o_lifm_l50)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(50), .NUMEL_LOG(6)
) vs_mt_50 (
    .i_vec(i_mt_l50), .stride(stride_l50), .o_vec(o_mt_l50)
);

// Shifter 51
wire [51*WORD_WIDTH-1:0] i_lifm_l51;
wire [51*WORD_WIDTH-1:0] o_lifm_l51;
wire [51*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l51;
wire [51*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l51;
wire [5:0] stride_l51;

assign i_lifm_l51 = {lifm_line_arr[50], 50*WORD_WIDTH'b0};
assign i_mt_l51 = {mt_line_arr[50], 50*WORD_WIDTH'b0};
assign stride_l51 = psum_arr[50][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(51), .NUMEL_LOG(6)
) vs_lifm_51 (
    .i_vec(i_lifm_l51), .stride(stride_l51), .o_vec(o_lifm_l51)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(51), .NUMEL_LOG(6)
) vs_mt_51 (
    .i_vec(i_mt_l51), .stride(stride_l51), .o_vec(o_mt_l51)
);

// Shifter 52
wire [52*WORD_WIDTH-1:0] i_lifm_l52;
wire [52*WORD_WIDTH-1:0] o_lifm_l52;
wire [52*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l52;
wire [52*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l52;
wire [5:0] stride_l52;

assign i_lifm_l52 = {lifm_line_arr[51], 51*WORD_WIDTH'b0};
assign i_mt_l52 = {mt_line_arr[51], 51*WORD_WIDTH'b0};
assign stride_l52 = psum_arr[51][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(52), .NUMEL_LOG(6)
) vs_lifm_52 (
    .i_vec(i_lifm_l52), .stride(stride_l52), .o_vec(o_lifm_l52)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(52), .NUMEL_LOG(6)
) vs_mt_52 (
    .i_vec(i_mt_l52), .stride(stride_l52), .o_vec(o_mt_l52)
);

// Shifter 53
wire [53*WORD_WIDTH-1:0] i_lifm_l53;
wire [53*WORD_WIDTH-1:0] o_lifm_l53;
wire [53*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l53;
wire [53*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l53;
wire [5:0] stride_l53;

assign i_lifm_l53 = {lifm_line_arr[52], 52*WORD_WIDTH'b0};
assign i_mt_l53 = {mt_line_arr[52], 52*WORD_WIDTH'b0};
assign stride_l53 = psum_arr[52][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(53), .NUMEL_LOG(6)
) vs_lifm_53 (
    .i_vec(i_lifm_l53), .stride(stride_l53), .o_vec(o_lifm_l53)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(53), .NUMEL_LOG(6)
) vs_mt_53 (
    .i_vec(i_mt_l53), .stride(stride_l53), .o_vec(o_mt_l53)
);

// Shifter 54
wire [54*WORD_WIDTH-1:0] i_lifm_l54;
wire [54*WORD_WIDTH-1:0] o_lifm_l54;
wire [54*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l54;
wire [54*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l54;
wire [5:0] stride_l54;

assign i_lifm_l54 = {lifm_line_arr[53], 53*WORD_WIDTH'b0};
assign i_mt_l54 = {mt_line_arr[53], 53*WORD_WIDTH'b0};
assign stride_l54 = psum_arr[53][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(54), .NUMEL_LOG(6)
) vs_lifm_54 (
    .i_vec(i_lifm_l54), .stride(stride_l54), .o_vec(o_lifm_l54)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(54), .NUMEL_LOG(6)
) vs_mt_54 (
    .i_vec(i_mt_l54), .stride(stride_l54), .o_vec(o_mt_l54)
);

// Shifter 55
wire [55*WORD_WIDTH-1:0] i_lifm_l55;
wire [55*WORD_WIDTH-1:0] o_lifm_l55;
wire [55*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l55;
wire [55*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l55;
wire [5:0] stride_l55;

assign i_lifm_l55 = {lifm_line_arr[54], 54*WORD_WIDTH'b0};
assign i_mt_l55 = {mt_line_arr[54], 54*WORD_WIDTH'b0};
assign stride_l55 = psum_arr[54][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(55), .NUMEL_LOG(6)
) vs_lifm_55 (
    .i_vec(i_lifm_l55), .stride(stride_l55), .o_vec(o_lifm_l55)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(55), .NUMEL_LOG(6)
) vs_mt_55 (
    .i_vec(i_mt_l55), .stride(stride_l55), .o_vec(o_mt_l55)
);

// Shifter 56
wire [56*WORD_WIDTH-1:0] i_lifm_l56;
wire [56*WORD_WIDTH-1:0] o_lifm_l56;
wire [56*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l56;
wire [56*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l56;
wire [5:0] stride_l56;

assign i_lifm_l56 = {lifm_line_arr[55], 55*WORD_WIDTH'b0};
assign i_mt_l56 = {mt_line_arr[55], 55*WORD_WIDTH'b0};
assign stride_l56 = psum_arr[55][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(56), .NUMEL_LOG(6)
) vs_lifm_56 (
    .i_vec(i_lifm_l56), .stride(stride_l56), .o_vec(o_lifm_l56)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(56), .NUMEL_LOG(6)
) vs_mt_56 (
    .i_vec(i_mt_l56), .stride(stride_l56), .o_vec(o_mt_l56)
);

// Shifter 57
wire [57*WORD_WIDTH-1:0] i_lifm_l57;
wire [57*WORD_WIDTH-1:0] o_lifm_l57;
wire [57*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l57;
wire [57*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l57;
wire [5:0] stride_l57;

assign i_lifm_l57 = {lifm_line_arr[56], 56*WORD_WIDTH'b0};
assign i_mt_l57 = {mt_line_arr[56], 56*WORD_WIDTH'b0};
assign stride_l57 = psum_arr[56][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(57), .NUMEL_LOG(6)
) vs_lifm_57 (
    .i_vec(i_lifm_l57), .stride(stride_l57), .o_vec(o_lifm_l57)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(57), .NUMEL_LOG(6)
) vs_mt_57 (
    .i_vec(i_mt_l57), .stride(stride_l57), .o_vec(o_mt_l57)
);

// Shifter 58
wire [58*WORD_WIDTH-1:0] i_lifm_l58;
wire [58*WORD_WIDTH-1:0] o_lifm_l58;
wire [58*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l58;
wire [58*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l58;
wire [5:0] stride_l58;

assign i_lifm_l58 = {lifm_line_arr[57], 57*WORD_WIDTH'b0};
assign i_mt_l58 = {mt_line_arr[57], 57*WORD_WIDTH'b0};
assign stride_l58 = psum_arr[57][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(58), .NUMEL_LOG(6)
) vs_lifm_58 (
    .i_vec(i_lifm_l58), .stride(stride_l58), .o_vec(o_lifm_l58)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(58), .NUMEL_LOG(6)
) vs_mt_58 (
    .i_vec(i_mt_l58), .stride(stride_l58), .o_vec(o_mt_l58)
);

// Shifter 59
wire [59*WORD_WIDTH-1:0] i_lifm_l59;
wire [59*WORD_WIDTH-1:0] o_lifm_l59;
wire [59*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l59;
wire [59*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l59;
wire [5:0] stride_l59;

assign i_lifm_l59 = {lifm_line_arr[58], 58*WORD_WIDTH'b0};
assign i_mt_l59 = {mt_line_arr[58], 58*WORD_WIDTH'b0};
assign stride_l59 = psum_arr[58][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(59), .NUMEL_LOG(6)
) vs_lifm_59 (
    .i_vec(i_lifm_l59), .stride(stride_l59), .o_vec(o_lifm_l59)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(59), .NUMEL_LOG(6)
) vs_mt_59 (
    .i_vec(i_mt_l59), .stride(stride_l59), .o_vec(o_mt_l59)
);

// Shifter 60
wire [60*WORD_WIDTH-1:0] i_lifm_l60;
wire [60*WORD_WIDTH-1:0] o_lifm_l60;
wire [60*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l60;
wire [60*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l60;
wire [5:0] stride_l60;

assign i_lifm_l60 = {lifm_line_arr[59], 59*WORD_WIDTH'b0};
assign i_mt_l60 = {mt_line_arr[59], 59*WORD_WIDTH'b0};
assign stride_l60 = psum_arr[59][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(60), .NUMEL_LOG(6)
) vs_lifm_60 (
    .i_vec(i_lifm_l60), .stride(stride_l60), .o_vec(o_lifm_l60)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(60), .NUMEL_LOG(6)
) vs_mt_60 (
    .i_vec(i_mt_l60), .stride(stride_l60), .o_vec(o_mt_l60)
);

// Shifter 61
wire [61*WORD_WIDTH-1:0] i_lifm_l61;
wire [61*WORD_WIDTH-1:0] o_lifm_l61;
wire [61*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l61;
wire [61*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l61;
wire [5:0] stride_l61;

assign i_lifm_l61 = {lifm_line_arr[60], 60*WORD_WIDTH'b0};
assign i_mt_l61 = {mt_line_arr[60], 60*WORD_WIDTH'b0};
assign stride_l61 = psum_arr[60][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(61), .NUMEL_LOG(6)
) vs_lifm_61 (
    .i_vec(i_lifm_l61), .stride(stride_l61), .o_vec(o_lifm_l61)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(61), .NUMEL_LOG(6)
) vs_mt_61 (
    .i_vec(i_mt_l61), .stride(stride_l61), .o_vec(o_mt_l61)
);

// Shifter 62
wire [62*WORD_WIDTH-1:0] i_lifm_l62;
wire [62*WORD_WIDTH-1:0] o_lifm_l62;
wire [62*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l62;
wire [62*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l62;
wire [5:0] stride_l62;

assign i_lifm_l62 = {lifm_line_arr[61], 61*WORD_WIDTH'b0};
assign i_mt_l62 = {mt_line_arr[61], 61*WORD_WIDTH'b0};
assign stride_l62 = psum_arr[61][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(62), .NUMEL_LOG(6)
) vs_lifm_62 (
    .i_vec(i_lifm_l62), .stride(stride_l62), .o_vec(o_lifm_l62)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(62), .NUMEL_LOG(6)
) vs_mt_62 (
    .i_vec(i_mt_l62), .stride(stride_l62), .o_vec(o_mt_l62)
);

// Shifter 63
wire [63*WORD_WIDTH-1:0] i_lifm_l63;
wire [63*WORD_WIDTH-1:0] o_lifm_l63;
wire [63*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l63;
wire [63*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l63;
wire [5:0] stride_l63;

assign i_lifm_l63 = {lifm_line_arr[62], 62*WORD_WIDTH'b0};
assign i_mt_l63 = {mt_line_arr[62], 62*WORD_WIDTH'b0};
assign stride_l63 = psum_arr[62][5:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(63), .NUMEL_LOG(6)
) vs_lifm_63 (
    .i_vec(i_lifm_l63), .stride(stride_l63), .o_vec(o_lifm_l63)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(63), .NUMEL_LOG(6)
) vs_mt_63 (
    .i_vec(i_mt_l63), .stride(stride_l63), .o_vec(o_mt_l63)
);

// Shifter 64
wire [64*WORD_WIDTH-1:0] i_lifm_l64;
wire [64*WORD_WIDTH-1:0] o_lifm_l64;
wire [64*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l64;
wire [64*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l64;
wire [6:0] stride_l64;

assign i_lifm_l64 = {lifm_line_arr[63], 63*WORD_WIDTH'b0};
assign i_mt_l64 = {mt_line_arr[63], 63*WORD_WIDTH'b0};
assign stride_l64 = psum_arr[63][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(64), .NUMEL_LOG(7)
) vs_lifm_64 (
    .i_vec(i_lifm_l64), .stride(stride_l64), .o_vec(o_lifm_l64)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(64), .NUMEL_LOG(7)
) vs_mt_64 (
    .i_vec(i_mt_l64), .stride(stride_l64), .o_vec(o_mt_l64)
);

// Shifter 65
wire [65*WORD_WIDTH-1:0] i_lifm_l65;
wire [65*WORD_WIDTH-1:0] o_lifm_l65;
wire [65*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l65;
wire [65*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l65;
wire [6:0] stride_l65;

assign i_lifm_l65 = {lifm_line_arr[64], 64*WORD_WIDTH'b0};
assign i_mt_l65 = {mt_line_arr[64], 64*WORD_WIDTH'b0};
assign stride_l65 = psum_arr[64][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(65), .NUMEL_LOG(7)
) vs_lifm_65 (
    .i_vec(i_lifm_l65), .stride(stride_l65), .o_vec(o_lifm_l65)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(65), .NUMEL_LOG(7)
) vs_mt_65 (
    .i_vec(i_mt_l65), .stride(stride_l65), .o_vec(o_mt_l65)
);

// Shifter 66
wire [66*WORD_WIDTH-1:0] i_lifm_l66;
wire [66*WORD_WIDTH-1:0] o_lifm_l66;
wire [66*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l66;
wire [66*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l66;
wire [6:0] stride_l66;

assign i_lifm_l66 = {lifm_line_arr[65], 65*WORD_WIDTH'b0};
assign i_mt_l66 = {mt_line_arr[65], 65*WORD_WIDTH'b0};
assign stride_l66 = psum_arr[65][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(66), .NUMEL_LOG(7)
) vs_lifm_66 (
    .i_vec(i_lifm_l66), .stride(stride_l66), .o_vec(o_lifm_l66)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(66), .NUMEL_LOG(7)
) vs_mt_66 (
    .i_vec(i_mt_l66), .stride(stride_l66), .o_vec(o_mt_l66)
);

// Shifter 67
wire [67*WORD_WIDTH-1:0] i_lifm_l67;
wire [67*WORD_WIDTH-1:0] o_lifm_l67;
wire [67*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l67;
wire [67*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l67;
wire [6:0] stride_l67;

assign i_lifm_l67 = {lifm_line_arr[66], 66*WORD_WIDTH'b0};
assign i_mt_l67 = {mt_line_arr[66], 66*WORD_WIDTH'b0};
assign stride_l67 = psum_arr[66][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(67), .NUMEL_LOG(7)
) vs_lifm_67 (
    .i_vec(i_lifm_l67), .stride(stride_l67), .o_vec(o_lifm_l67)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(67), .NUMEL_LOG(7)
) vs_mt_67 (
    .i_vec(i_mt_l67), .stride(stride_l67), .o_vec(o_mt_l67)
);

// Shifter 68
wire [68*WORD_WIDTH-1:0] i_lifm_l68;
wire [68*WORD_WIDTH-1:0] o_lifm_l68;
wire [68*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l68;
wire [68*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l68;
wire [6:0] stride_l68;

assign i_lifm_l68 = {lifm_line_arr[67], 67*WORD_WIDTH'b0};
assign i_mt_l68 = {mt_line_arr[67], 67*WORD_WIDTH'b0};
assign stride_l68 = psum_arr[67][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(68), .NUMEL_LOG(7)
) vs_lifm_68 (
    .i_vec(i_lifm_l68), .stride(stride_l68), .o_vec(o_lifm_l68)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(68), .NUMEL_LOG(7)
) vs_mt_68 (
    .i_vec(i_mt_l68), .stride(stride_l68), .o_vec(o_mt_l68)
);

// Shifter 69
wire [69*WORD_WIDTH-1:0] i_lifm_l69;
wire [69*WORD_WIDTH-1:0] o_lifm_l69;
wire [69*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l69;
wire [69*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l69;
wire [6:0] stride_l69;

assign i_lifm_l69 = {lifm_line_arr[68], 68*WORD_WIDTH'b0};
assign i_mt_l69 = {mt_line_arr[68], 68*WORD_WIDTH'b0};
assign stride_l69 = psum_arr[68][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(69), .NUMEL_LOG(7)
) vs_lifm_69 (
    .i_vec(i_lifm_l69), .stride(stride_l69), .o_vec(o_lifm_l69)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(69), .NUMEL_LOG(7)
) vs_mt_69 (
    .i_vec(i_mt_l69), .stride(stride_l69), .o_vec(o_mt_l69)
);

// Shifter 70
wire [70*WORD_WIDTH-1:0] i_lifm_l70;
wire [70*WORD_WIDTH-1:0] o_lifm_l70;
wire [70*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l70;
wire [70*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l70;
wire [6:0] stride_l70;

assign i_lifm_l70 = {lifm_line_arr[69], 69*WORD_WIDTH'b0};
assign i_mt_l70 = {mt_line_arr[69], 69*WORD_WIDTH'b0};
assign stride_l70 = psum_arr[69][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(70), .NUMEL_LOG(7)
) vs_lifm_70 (
    .i_vec(i_lifm_l70), .stride(stride_l70), .o_vec(o_lifm_l70)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(70), .NUMEL_LOG(7)
) vs_mt_70 (
    .i_vec(i_mt_l70), .stride(stride_l70), .o_vec(o_mt_l70)
);

// Shifter 71
wire [71*WORD_WIDTH-1:0] i_lifm_l71;
wire [71*WORD_WIDTH-1:0] o_lifm_l71;
wire [71*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l71;
wire [71*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l71;
wire [6:0] stride_l71;

assign i_lifm_l71 = {lifm_line_arr[70], 70*WORD_WIDTH'b0};
assign i_mt_l71 = {mt_line_arr[70], 70*WORD_WIDTH'b0};
assign stride_l71 = psum_arr[70][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(71), .NUMEL_LOG(7)
) vs_lifm_71 (
    .i_vec(i_lifm_l71), .stride(stride_l71), .o_vec(o_lifm_l71)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(71), .NUMEL_LOG(7)
) vs_mt_71 (
    .i_vec(i_mt_l71), .stride(stride_l71), .o_vec(o_mt_l71)
);

// Shifter 72
wire [72*WORD_WIDTH-1:0] i_lifm_l72;
wire [72*WORD_WIDTH-1:0] o_lifm_l72;
wire [72*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l72;
wire [72*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l72;
wire [6:0] stride_l72;

assign i_lifm_l72 = {lifm_line_arr[71], 71*WORD_WIDTH'b0};
assign i_mt_l72 = {mt_line_arr[71], 71*WORD_WIDTH'b0};
assign stride_l72 = psum_arr[71][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(72), .NUMEL_LOG(7)
) vs_lifm_72 (
    .i_vec(i_lifm_l72), .stride(stride_l72), .o_vec(o_lifm_l72)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(72), .NUMEL_LOG(7)
) vs_mt_72 (
    .i_vec(i_mt_l72), .stride(stride_l72), .o_vec(o_mt_l72)
);

// Shifter 73
wire [73*WORD_WIDTH-1:0] i_lifm_l73;
wire [73*WORD_WIDTH-1:0] o_lifm_l73;
wire [73*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l73;
wire [73*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l73;
wire [6:0] stride_l73;

assign i_lifm_l73 = {lifm_line_arr[72], 72*WORD_WIDTH'b0};
assign i_mt_l73 = {mt_line_arr[72], 72*WORD_WIDTH'b0};
assign stride_l73 = psum_arr[72][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(73), .NUMEL_LOG(7)
) vs_lifm_73 (
    .i_vec(i_lifm_l73), .stride(stride_l73), .o_vec(o_lifm_l73)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(73), .NUMEL_LOG(7)
) vs_mt_73 (
    .i_vec(i_mt_l73), .stride(stride_l73), .o_vec(o_mt_l73)
);

// Shifter 74
wire [74*WORD_WIDTH-1:0] i_lifm_l74;
wire [74*WORD_WIDTH-1:0] o_lifm_l74;
wire [74*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l74;
wire [74*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l74;
wire [6:0] stride_l74;

assign i_lifm_l74 = {lifm_line_arr[73], 73*WORD_WIDTH'b0};
assign i_mt_l74 = {mt_line_arr[73], 73*WORD_WIDTH'b0};
assign stride_l74 = psum_arr[73][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(74), .NUMEL_LOG(7)
) vs_lifm_74 (
    .i_vec(i_lifm_l74), .stride(stride_l74), .o_vec(o_lifm_l74)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(74), .NUMEL_LOG(7)
) vs_mt_74 (
    .i_vec(i_mt_l74), .stride(stride_l74), .o_vec(o_mt_l74)
);

// Shifter 75
wire [75*WORD_WIDTH-1:0] i_lifm_l75;
wire [75*WORD_WIDTH-1:0] o_lifm_l75;
wire [75*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l75;
wire [75*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l75;
wire [6:0] stride_l75;

assign i_lifm_l75 = {lifm_line_arr[74], 74*WORD_WIDTH'b0};
assign i_mt_l75 = {mt_line_arr[74], 74*WORD_WIDTH'b0};
assign stride_l75 = psum_arr[74][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(75), .NUMEL_LOG(7)
) vs_lifm_75 (
    .i_vec(i_lifm_l75), .stride(stride_l75), .o_vec(o_lifm_l75)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(75), .NUMEL_LOG(7)
) vs_mt_75 (
    .i_vec(i_mt_l75), .stride(stride_l75), .o_vec(o_mt_l75)
);

// Shifter 76
wire [76*WORD_WIDTH-1:0] i_lifm_l76;
wire [76*WORD_WIDTH-1:0] o_lifm_l76;
wire [76*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l76;
wire [76*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l76;
wire [6:0] stride_l76;

assign i_lifm_l76 = {lifm_line_arr[75], 75*WORD_WIDTH'b0};
assign i_mt_l76 = {mt_line_arr[75], 75*WORD_WIDTH'b0};
assign stride_l76 = psum_arr[75][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(76), .NUMEL_LOG(7)
) vs_lifm_76 (
    .i_vec(i_lifm_l76), .stride(stride_l76), .o_vec(o_lifm_l76)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(76), .NUMEL_LOG(7)
) vs_mt_76 (
    .i_vec(i_mt_l76), .stride(stride_l76), .o_vec(o_mt_l76)
);

// Shifter 77
wire [77*WORD_WIDTH-1:0] i_lifm_l77;
wire [77*WORD_WIDTH-1:0] o_lifm_l77;
wire [77*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l77;
wire [77*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l77;
wire [6:0] stride_l77;

assign i_lifm_l77 = {lifm_line_arr[76], 76*WORD_WIDTH'b0};
assign i_mt_l77 = {mt_line_arr[76], 76*WORD_WIDTH'b0};
assign stride_l77 = psum_arr[76][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(77), .NUMEL_LOG(7)
) vs_lifm_77 (
    .i_vec(i_lifm_l77), .stride(stride_l77), .o_vec(o_lifm_l77)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(77), .NUMEL_LOG(7)
) vs_mt_77 (
    .i_vec(i_mt_l77), .stride(stride_l77), .o_vec(o_mt_l77)
);

// Shifter 78
wire [78*WORD_WIDTH-1:0] i_lifm_l78;
wire [78*WORD_WIDTH-1:0] o_lifm_l78;
wire [78*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l78;
wire [78*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l78;
wire [6:0] stride_l78;

assign i_lifm_l78 = {lifm_line_arr[77], 77*WORD_WIDTH'b0};
assign i_mt_l78 = {mt_line_arr[77], 77*WORD_WIDTH'b0};
assign stride_l78 = psum_arr[77][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(78), .NUMEL_LOG(7)
) vs_lifm_78 (
    .i_vec(i_lifm_l78), .stride(stride_l78), .o_vec(o_lifm_l78)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(78), .NUMEL_LOG(7)
) vs_mt_78 (
    .i_vec(i_mt_l78), .stride(stride_l78), .o_vec(o_mt_l78)
);

// Shifter 79
wire [79*WORD_WIDTH-1:0] i_lifm_l79;
wire [79*WORD_WIDTH-1:0] o_lifm_l79;
wire [79*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l79;
wire [79*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l79;
wire [6:0] stride_l79;

assign i_lifm_l79 = {lifm_line_arr[78], 78*WORD_WIDTH'b0};
assign i_mt_l79 = {mt_line_arr[78], 78*WORD_WIDTH'b0};
assign stride_l79 = psum_arr[78][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(79), .NUMEL_LOG(7)
) vs_lifm_79 (
    .i_vec(i_lifm_l79), .stride(stride_l79), .o_vec(o_lifm_l79)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(79), .NUMEL_LOG(7)
) vs_mt_79 (
    .i_vec(i_mt_l79), .stride(stride_l79), .o_vec(o_mt_l79)
);

// Shifter 80
wire [80*WORD_WIDTH-1:0] i_lifm_l80;
wire [80*WORD_WIDTH-1:0] o_lifm_l80;
wire [80*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l80;
wire [80*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l80;
wire [6:0] stride_l80;

assign i_lifm_l80 = {lifm_line_arr[79], 79*WORD_WIDTH'b0};
assign i_mt_l80 = {mt_line_arr[79], 79*WORD_WIDTH'b0};
assign stride_l80 = psum_arr[79][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(80), .NUMEL_LOG(7)
) vs_lifm_80 (
    .i_vec(i_lifm_l80), .stride(stride_l80), .o_vec(o_lifm_l80)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(80), .NUMEL_LOG(7)
) vs_mt_80 (
    .i_vec(i_mt_l80), .stride(stride_l80), .o_vec(o_mt_l80)
);

// Shifter 81
wire [81*WORD_WIDTH-1:0] i_lifm_l81;
wire [81*WORD_WIDTH-1:0] o_lifm_l81;
wire [81*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l81;
wire [81*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l81;
wire [6:0] stride_l81;

assign i_lifm_l81 = {lifm_line_arr[80], 80*WORD_WIDTH'b0};
assign i_mt_l81 = {mt_line_arr[80], 80*WORD_WIDTH'b0};
assign stride_l81 = psum_arr[80][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(81), .NUMEL_LOG(7)
) vs_lifm_81 (
    .i_vec(i_lifm_l81), .stride(stride_l81), .o_vec(o_lifm_l81)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(81), .NUMEL_LOG(7)
) vs_mt_81 (
    .i_vec(i_mt_l81), .stride(stride_l81), .o_vec(o_mt_l81)
);

// Shifter 82
wire [82*WORD_WIDTH-1:0] i_lifm_l82;
wire [82*WORD_WIDTH-1:0] o_lifm_l82;
wire [82*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l82;
wire [82*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l82;
wire [6:0] stride_l82;

assign i_lifm_l82 = {lifm_line_arr[81], 81*WORD_WIDTH'b0};
assign i_mt_l82 = {mt_line_arr[81], 81*WORD_WIDTH'b0};
assign stride_l82 = psum_arr[81][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(82), .NUMEL_LOG(7)
) vs_lifm_82 (
    .i_vec(i_lifm_l82), .stride(stride_l82), .o_vec(o_lifm_l82)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(82), .NUMEL_LOG(7)
) vs_mt_82 (
    .i_vec(i_mt_l82), .stride(stride_l82), .o_vec(o_mt_l82)
);

// Shifter 83
wire [83*WORD_WIDTH-1:0] i_lifm_l83;
wire [83*WORD_WIDTH-1:0] o_lifm_l83;
wire [83*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l83;
wire [83*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l83;
wire [6:0] stride_l83;

assign i_lifm_l83 = {lifm_line_arr[82], 82*WORD_WIDTH'b0};
assign i_mt_l83 = {mt_line_arr[82], 82*WORD_WIDTH'b0};
assign stride_l83 = psum_arr[82][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(83), .NUMEL_LOG(7)
) vs_lifm_83 (
    .i_vec(i_lifm_l83), .stride(stride_l83), .o_vec(o_lifm_l83)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(83), .NUMEL_LOG(7)
) vs_mt_83 (
    .i_vec(i_mt_l83), .stride(stride_l83), .o_vec(o_mt_l83)
);

// Shifter 84
wire [84*WORD_WIDTH-1:0] i_lifm_l84;
wire [84*WORD_WIDTH-1:0] o_lifm_l84;
wire [84*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l84;
wire [84*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l84;
wire [6:0] stride_l84;

assign i_lifm_l84 = {lifm_line_arr[83], 83*WORD_WIDTH'b0};
assign i_mt_l84 = {mt_line_arr[83], 83*WORD_WIDTH'b0};
assign stride_l84 = psum_arr[83][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(84), .NUMEL_LOG(7)
) vs_lifm_84 (
    .i_vec(i_lifm_l84), .stride(stride_l84), .o_vec(o_lifm_l84)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(84), .NUMEL_LOG(7)
) vs_mt_84 (
    .i_vec(i_mt_l84), .stride(stride_l84), .o_vec(o_mt_l84)
);

// Shifter 85
wire [85*WORD_WIDTH-1:0] i_lifm_l85;
wire [85*WORD_WIDTH-1:0] o_lifm_l85;
wire [85*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l85;
wire [85*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l85;
wire [6:0] stride_l85;

assign i_lifm_l85 = {lifm_line_arr[84], 84*WORD_WIDTH'b0};
assign i_mt_l85 = {mt_line_arr[84], 84*WORD_WIDTH'b0};
assign stride_l85 = psum_arr[84][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(85), .NUMEL_LOG(7)
) vs_lifm_85 (
    .i_vec(i_lifm_l85), .stride(stride_l85), .o_vec(o_lifm_l85)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(85), .NUMEL_LOG(7)
) vs_mt_85 (
    .i_vec(i_mt_l85), .stride(stride_l85), .o_vec(o_mt_l85)
);

// Shifter 86
wire [86*WORD_WIDTH-1:0] i_lifm_l86;
wire [86*WORD_WIDTH-1:0] o_lifm_l86;
wire [86*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l86;
wire [86*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l86;
wire [6:0] stride_l86;

assign i_lifm_l86 = {lifm_line_arr[85], 85*WORD_WIDTH'b0};
assign i_mt_l86 = {mt_line_arr[85], 85*WORD_WIDTH'b0};
assign stride_l86 = psum_arr[85][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(86), .NUMEL_LOG(7)
) vs_lifm_86 (
    .i_vec(i_lifm_l86), .stride(stride_l86), .o_vec(o_lifm_l86)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(86), .NUMEL_LOG(7)
) vs_mt_86 (
    .i_vec(i_mt_l86), .stride(stride_l86), .o_vec(o_mt_l86)
);

// Shifter 87
wire [87*WORD_WIDTH-1:0] i_lifm_l87;
wire [87*WORD_WIDTH-1:0] o_lifm_l87;
wire [87*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l87;
wire [87*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l87;
wire [6:0] stride_l87;

assign i_lifm_l87 = {lifm_line_arr[86], 86*WORD_WIDTH'b0};
assign i_mt_l87 = {mt_line_arr[86], 86*WORD_WIDTH'b0};
assign stride_l87 = psum_arr[86][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(87), .NUMEL_LOG(7)
) vs_lifm_87 (
    .i_vec(i_lifm_l87), .stride(stride_l87), .o_vec(o_lifm_l87)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(87), .NUMEL_LOG(7)
) vs_mt_87 (
    .i_vec(i_mt_l87), .stride(stride_l87), .o_vec(o_mt_l87)
);

// Shifter 88
wire [88*WORD_WIDTH-1:0] i_lifm_l88;
wire [88*WORD_WIDTH-1:0] o_lifm_l88;
wire [88*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l88;
wire [88*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l88;
wire [6:0] stride_l88;

assign i_lifm_l88 = {lifm_line_arr[87], 87*WORD_WIDTH'b0};
assign i_mt_l88 = {mt_line_arr[87], 87*WORD_WIDTH'b0};
assign stride_l88 = psum_arr[87][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(88), .NUMEL_LOG(7)
) vs_lifm_88 (
    .i_vec(i_lifm_l88), .stride(stride_l88), .o_vec(o_lifm_l88)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(88), .NUMEL_LOG(7)
) vs_mt_88 (
    .i_vec(i_mt_l88), .stride(stride_l88), .o_vec(o_mt_l88)
);

// Shifter 89
wire [89*WORD_WIDTH-1:0] i_lifm_l89;
wire [89*WORD_WIDTH-1:0] o_lifm_l89;
wire [89*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l89;
wire [89*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l89;
wire [6:0] stride_l89;

assign i_lifm_l89 = {lifm_line_arr[88], 88*WORD_WIDTH'b0};
assign i_mt_l89 = {mt_line_arr[88], 88*WORD_WIDTH'b0};
assign stride_l89 = psum_arr[88][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(89), .NUMEL_LOG(7)
) vs_lifm_89 (
    .i_vec(i_lifm_l89), .stride(stride_l89), .o_vec(o_lifm_l89)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(89), .NUMEL_LOG(7)
) vs_mt_89 (
    .i_vec(i_mt_l89), .stride(stride_l89), .o_vec(o_mt_l89)
);

// Shifter 90
wire [90*WORD_WIDTH-1:0] i_lifm_l90;
wire [90*WORD_WIDTH-1:0] o_lifm_l90;
wire [90*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l90;
wire [90*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l90;
wire [6:0] stride_l90;

assign i_lifm_l90 = {lifm_line_arr[89], 89*WORD_WIDTH'b0};
assign i_mt_l90 = {mt_line_arr[89], 89*WORD_WIDTH'b0};
assign stride_l90 = psum_arr[89][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(90), .NUMEL_LOG(7)
) vs_lifm_90 (
    .i_vec(i_lifm_l90), .stride(stride_l90), .o_vec(o_lifm_l90)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(90), .NUMEL_LOG(7)
) vs_mt_90 (
    .i_vec(i_mt_l90), .stride(stride_l90), .o_vec(o_mt_l90)
);

// Shifter 91
wire [91*WORD_WIDTH-1:0] i_lifm_l91;
wire [91*WORD_WIDTH-1:0] o_lifm_l91;
wire [91*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l91;
wire [91*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l91;
wire [6:0] stride_l91;

assign i_lifm_l91 = {lifm_line_arr[90], 90*WORD_WIDTH'b0};
assign i_mt_l91 = {mt_line_arr[90], 90*WORD_WIDTH'b0};
assign stride_l91 = psum_arr[90][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(91), .NUMEL_LOG(7)
) vs_lifm_91 (
    .i_vec(i_lifm_l91), .stride(stride_l91), .o_vec(o_lifm_l91)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(91), .NUMEL_LOG(7)
) vs_mt_91 (
    .i_vec(i_mt_l91), .stride(stride_l91), .o_vec(o_mt_l91)
);

// Shifter 92
wire [92*WORD_WIDTH-1:0] i_lifm_l92;
wire [92*WORD_WIDTH-1:0] o_lifm_l92;
wire [92*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l92;
wire [92*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l92;
wire [6:0] stride_l92;

assign i_lifm_l92 = {lifm_line_arr[91], 91*WORD_WIDTH'b0};
assign i_mt_l92 = {mt_line_arr[91], 91*WORD_WIDTH'b0};
assign stride_l92 = psum_arr[91][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(92), .NUMEL_LOG(7)
) vs_lifm_92 (
    .i_vec(i_lifm_l92), .stride(stride_l92), .o_vec(o_lifm_l92)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(92), .NUMEL_LOG(7)
) vs_mt_92 (
    .i_vec(i_mt_l92), .stride(stride_l92), .o_vec(o_mt_l92)
);

// Shifter 93
wire [93*WORD_WIDTH-1:0] i_lifm_l93;
wire [93*WORD_WIDTH-1:0] o_lifm_l93;
wire [93*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l93;
wire [93*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l93;
wire [6:0] stride_l93;

assign i_lifm_l93 = {lifm_line_arr[92], 92*WORD_WIDTH'b0};
assign i_mt_l93 = {mt_line_arr[92], 92*WORD_WIDTH'b0};
assign stride_l93 = psum_arr[92][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(93), .NUMEL_LOG(7)
) vs_lifm_93 (
    .i_vec(i_lifm_l93), .stride(stride_l93), .o_vec(o_lifm_l93)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(93), .NUMEL_LOG(7)
) vs_mt_93 (
    .i_vec(i_mt_l93), .stride(stride_l93), .o_vec(o_mt_l93)
);

// Shifter 94
wire [94*WORD_WIDTH-1:0] i_lifm_l94;
wire [94*WORD_WIDTH-1:0] o_lifm_l94;
wire [94*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l94;
wire [94*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l94;
wire [6:0] stride_l94;

assign i_lifm_l94 = {lifm_line_arr[93], 93*WORD_WIDTH'b0};
assign i_mt_l94 = {mt_line_arr[93], 93*WORD_WIDTH'b0};
assign stride_l94 = psum_arr[93][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(94), .NUMEL_LOG(7)
) vs_lifm_94 (
    .i_vec(i_lifm_l94), .stride(stride_l94), .o_vec(o_lifm_l94)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(94), .NUMEL_LOG(7)
) vs_mt_94 (
    .i_vec(i_mt_l94), .stride(stride_l94), .o_vec(o_mt_l94)
);

// Shifter 95
wire [95*WORD_WIDTH-1:0] i_lifm_l95;
wire [95*WORD_WIDTH-1:0] o_lifm_l95;
wire [95*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l95;
wire [95*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l95;
wire [6:0] stride_l95;

assign i_lifm_l95 = {lifm_line_arr[94], 94*WORD_WIDTH'b0};
assign i_mt_l95 = {mt_line_arr[94], 94*WORD_WIDTH'b0};
assign stride_l95 = psum_arr[94][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(95), .NUMEL_LOG(7)
) vs_lifm_95 (
    .i_vec(i_lifm_l95), .stride(stride_l95), .o_vec(o_lifm_l95)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(95), .NUMEL_LOG(7)
) vs_mt_95 (
    .i_vec(i_mt_l95), .stride(stride_l95), .o_vec(o_mt_l95)
);

// Shifter 96
wire [96*WORD_WIDTH-1:0] i_lifm_l96;
wire [96*WORD_WIDTH-1:0] o_lifm_l96;
wire [96*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l96;
wire [96*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l96;
wire [6:0] stride_l96;

assign i_lifm_l96 = {lifm_line_arr[95], 95*WORD_WIDTH'b0};
assign i_mt_l96 = {mt_line_arr[95], 95*WORD_WIDTH'b0};
assign stride_l96 = psum_arr[95][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(96), .NUMEL_LOG(7)
) vs_lifm_96 (
    .i_vec(i_lifm_l96), .stride(stride_l96), .o_vec(o_lifm_l96)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(96), .NUMEL_LOG(7)
) vs_mt_96 (
    .i_vec(i_mt_l96), .stride(stride_l96), .o_vec(o_mt_l96)
);

// Shifter 97
wire [97*WORD_WIDTH-1:0] i_lifm_l97;
wire [97*WORD_WIDTH-1:0] o_lifm_l97;
wire [97*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l97;
wire [97*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l97;
wire [6:0] stride_l97;

assign i_lifm_l97 = {lifm_line_arr[96], 96*WORD_WIDTH'b0};
assign i_mt_l97 = {mt_line_arr[96], 96*WORD_WIDTH'b0};
assign stride_l97 = psum_arr[96][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(97), .NUMEL_LOG(7)
) vs_lifm_97 (
    .i_vec(i_lifm_l97), .stride(stride_l97), .o_vec(o_lifm_l97)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(97), .NUMEL_LOG(7)
) vs_mt_97 (
    .i_vec(i_mt_l97), .stride(stride_l97), .o_vec(o_mt_l97)
);

// Shifter 98
wire [98*WORD_WIDTH-1:0] i_lifm_l98;
wire [98*WORD_WIDTH-1:0] o_lifm_l98;
wire [98*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l98;
wire [98*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l98;
wire [6:0] stride_l98;

assign i_lifm_l98 = {lifm_line_arr[97], 97*WORD_WIDTH'b0};
assign i_mt_l98 = {mt_line_arr[97], 97*WORD_WIDTH'b0};
assign stride_l98 = psum_arr[97][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(98), .NUMEL_LOG(7)
) vs_lifm_98 (
    .i_vec(i_lifm_l98), .stride(stride_l98), .o_vec(o_lifm_l98)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(98), .NUMEL_LOG(7)
) vs_mt_98 (
    .i_vec(i_mt_l98), .stride(stride_l98), .o_vec(o_mt_l98)
);

// Shifter 99
wire [99*WORD_WIDTH-1:0] i_lifm_l99;
wire [99*WORD_WIDTH-1:0] o_lifm_l99;
wire [99*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l99;
wire [99*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l99;
wire [6:0] stride_l99;

assign i_lifm_l99 = {lifm_line_arr[98], 98*WORD_WIDTH'b0};
assign i_mt_l99 = {mt_line_arr[98], 98*WORD_WIDTH'b0};
assign stride_l99 = psum_arr[98][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(99), .NUMEL_LOG(7)
) vs_lifm_99 (
    .i_vec(i_lifm_l99), .stride(stride_l99), .o_vec(o_lifm_l99)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(99), .NUMEL_LOG(7)
) vs_mt_99 (
    .i_vec(i_mt_l99), .stride(stride_l99), .o_vec(o_mt_l99)
);

// Shifter 100
wire [100*WORD_WIDTH-1:0] i_lifm_l100;
wire [100*WORD_WIDTH-1:0] o_lifm_l100;
wire [100*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l100;
wire [100*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l100;
wire [6:0] stride_l100;

assign i_lifm_l100 = {lifm_line_arr[99], 99*WORD_WIDTH'b0};
assign i_mt_l100 = {mt_line_arr[99], 99*WORD_WIDTH'b0};
assign stride_l100 = psum_arr[99][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(100), .NUMEL_LOG(7)
) vs_lifm_100 (
    .i_vec(i_lifm_l100), .stride(stride_l100), .o_vec(o_lifm_l100)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(100), .NUMEL_LOG(7)
) vs_mt_100 (
    .i_vec(i_mt_l100), .stride(stride_l100), .o_vec(o_mt_l100)
);

// Shifter 101
wire [101*WORD_WIDTH-1:0] i_lifm_l101;
wire [101*WORD_WIDTH-1:0] o_lifm_l101;
wire [101*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l101;
wire [101*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l101;
wire [6:0] stride_l101;

assign i_lifm_l101 = {lifm_line_arr[100], 100*WORD_WIDTH'b0};
assign i_mt_l101 = {mt_line_arr[100], 100*WORD_WIDTH'b0};
assign stride_l101 = psum_arr[100][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(101), .NUMEL_LOG(7)
) vs_lifm_101 (
    .i_vec(i_lifm_l101), .stride(stride_l101), .o_vec(o_lifm_l101)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(101), .NUMEL_LOG(7)
) vs_mt_101 (
    .i_vec(i_mt_l101), .stride(stride_l101), .o_vec(o_mt_l101)
);

// Shifter 102
wire [102*WORD_WIDTH-1:0] i_lifm_l102;
wire [102*WORD_WIDTH-1:0] o_lifm_l102;
wire [102*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l102;
wire [102*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l102;
wire [6:0] stride_l102;

assign i_lifm_l102 = {lifm_line_arr[101], 101*WORD_WIDTH'b0};
assign i_mt_l102 = {mt_line_arr[101], 101*WORD_WIDTH'b0};
assign stride_l102 = psum_arr[101][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(102), .NUMEL_LOG(7)
) vs_lifm_102 (
    .i_vec(i_lifm_l102), .stride(stride_l102), .o_vec(o_lifm_l102)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(102), .NUMEL_LOG(7)
) vs_mt_102 (
    .i_vec(i_mt_l102), .stride(stride_l102), .o_vec(o_mt_l102)
);

// Shifter 103
wire [103*WORD_WIDTH-1:0] i_lifm_l103;
wire [103*WORD_WIDTH-1:0] o_lifm_l103;
wire [103*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l103;
wire [103*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l103;
wire [6:0] stride_l103;

assign i_lifm_l103 = {lifm_line_arr[102], 102*WORD_WIDTH'b0};
assign i_mt_l103 = {mt_line_arr[102], 102*WORD_WIDTH'b0};
assign stride_l103 = psum_arr[102][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(103), .NUMEL_LOG(7)
) vs_lifm_103 (
    .i_vec(i_lifm_l103), .stride(stride_l103), .o_vec(o_lifm_l103)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(103), .NUMEL_LOG(7)
) vs_mt_103 (
    .i_vec(i_mt_l103), .stride(stride_l103), .o_vec(o_mt_l103)
);

// Shifter 104
wire [104*WORD_WIDTH-1:0] i_lifm_l104;
wire [104*WORD_WIDTH-1:0] o_lifm_l104;
wire [104*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l104;
wire [104*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l104;
wire [6:0] stride_l104;

assign i_lifm_l104 = {lifm_line_arr[103], 103*WORD_WIDTH'b0};
assign i_mt_l104 = {mt_line_arr[103], 103*WORD_WIDTH'b0};
assign stride_l104 = psum_arr[103][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(104), .NUMEL_LOG(7)
) vs_lifm_104 (
    .i_vec(i_lifm_l104), .stride(stride_l104), .o_vec(o_lifm_l104)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(104), .NUMEL_LOG(7)
) vs_mt_104 (
    .i_vec(i_mt_l104), .stride(stride_l104), .o_vec(o_mt_l104)
);

// Shifter 105
wire [105*WORD_WIDTH-1:0] i_lifm_l105;
wire [105*WORD_WIDTH-1:0] o_lifm_l105;
wire [105*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l105;
wire [105*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l105;
wire [6:0] stride_l105;

assign i_lifm_l105 = {lifm_line_arr[104], 104*WORD_WIDTH'b0};
assign i_mt_l105 = {mt_line_arr[104], 104*WORD_WIDTH'b0};
assign stride_l105 = psum_arr[104][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(105), .NUMEL_LOG(7)
) vs_lifm_105 (
    .i_vec(i_lifm_l105), .stride(stride_l105), .o_vec(o_lifm_l105)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(105), .NUMEL_LOG(7)
) vs_mt_105 (
    .i_vec(i_mt_l105), .stride(stride_l105), .o_vec(o_mt_l105)
);

// Shifter 106
wire [106*WORD_WIDTH-1:0] i_lifm_l106;
wire [106*WORD_WIDTH-1:0] o_lifm_l106;
wire [106*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l106;
wire [106*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l106;
wire [6:0] stride_l106;

assign i_lifm_l106 = {lifm_line_arr[105], 105*WORD_WIDTH'b0};
assign i_mt_l106 = {mt_line_arr[105], 105*WORD_WIDTH'b0};
assign stride_l106 = psum_arr[105][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(106), .NUMEL_LOG(7)
) vs_lifm_106 (
    .i_vec(i_lifm_l106), .stride(stride_l106), .o_vec(o_lifm_l106)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(106), .NUMEL_LOG(7)
) vs_mt_106 (
    .i_vec(i_mt_l106), .stride(stride_l106), .o_vec(o_mt_l106)
);

// Shifter 107
wire [107*WORD_WIDTH-1:0] i_lifm_l107;
wire [107*WORD_WIDTH-1:0] o_lifm_l107;
wire [107*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l107;
wire [107*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l107;
wire [6:0] stride_l107;

assign i_lifm_l107 = {lifm_line_arr[106], 106*WORD_WIDTH'b0};
assign i_mt_l107 = {mt_line_arr[106], 106*WORD_WIDTH'b0};
assign stride_l107 = psum_arr[106][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(107), .NUMEL_LOG(7)
) vs_lifm_107 (
    .i_vec(i_lifm_l107), .stride(stride_l107), .o_vec(o_lifm_l107)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(107), .NUMEL_LOG(7)
) vs_mt_107 (
    .i_vec(i_mt_l107), .stride(stride_l107), .o_vec(o_mt_l107)
);

// Shifter 108
wire [108*WORD_WIDTH-1:0] i_lifm_l108;
wire [108*WORD_WIDTH-1:0] o_lifm_l108;
wire [108*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l108;
wire [108*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l108;
wire [6:0] stride_l108;

assign i_lifm_l108 = {lifm_line_arr[107], 107*WORD_WIDTH'b0};
assign i_mt_l108 = {mt_line_arr[107], 107*WORD_WIDTH'b0};
assign stride_l108 = psum_arr[107][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(108), .NUMEL_LOG(7)
) vs_lifm_108 (
    .i_vec(i_lifm_l108), .stride(stride_l108), .o_vec(o_lifm_l108)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(108), .NUMEL_LOG(7)
) vs_mt_108 (
    .i_vec(i_mt_l108), .stride(stride_l108), .o_vec(o_mt_l108)
);

// Shifter 109
wire [109*WORD_WIDTH-1:0] i_lifm_l109;
wire [109*WORD_WIDTH-1:0] o_lifm_l109;
wire [109*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l109;
wire [109*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l109;
wire [6:0] stride_l109;

assign i_lifm_l109 = {lifm_line_arr[108], 108*WORD_WIDTH'b0};
assign i_mt_l109 = {mt_line_arr[108], 108*WORD_WIDTH'b0};
assign stride_l109 = psum_arr[108][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(109), .NUMEL_LOG(7)
) vs_lifm_109 (
    .i_vec(i_lifm_l109), .stride(stride_l109), .o_vec(o_lifm_l109)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(109), .NUMEL_LOG(7)
) vs_mt_109 (
    .i_vec(i_mt_l109), .stride(stride_l109), .o_vec(o_mt_l109)
);

// Shifter 110
wire [110*WORD_WIDTH-1:0] i_lifm_l110;
wire [110*WORD_WIDTH-1:0] o_lifm_l110;
wire [110*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l110;
wire [110*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l110;
wire [6:0] stride_l110;

assign i_lifm_l110 = {lifm_line_arr[109], 109*WORD_WIDTH'b0};
assign i_mt_l110 = {mt_line_arr[109], 109*WORD_WIDTH'b0};
assign stride_l110 = psum_arr[109][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(110), .NUMEL_LOG(7)
) vs_lifm_110 (
    .i_vec(i_lifm_l110), .stride(stride_l110), .o_vec(o_lifm_l110)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(110), .NUMEL_LOG(7)
) vs_mt_110 (
    .i_vec(i_mt_l110), .stride(stride_l110), .o_vec(o_mt_l110)
);

// Shifter 111
wire [111*WORD_WIDTH-1:0] i_lifm_l111;
wire [111*WORD_WIDTH-1:0] o_lifm_l111;
wire [111*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l111;
wire [111*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l111;
wire [6:0] stride_l111;

assign i_lifm_l111 = {lifm_line_arr[110], 110*WORD_WIDTH'b0};
assign i_mt_l111 = {mt_line_arr[110], 110*WORD_WIDTH'b0};
assign stride_l111 = psum_arr[110][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(111), .NUMEL_LOG(7)
) vs_lifm_111 (
    .i_vec(i_lifm_l111), .stride(stride_l111), .o_vec(o_lifm_l111)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(111), .NUMEL_LOG(7)
) vs_mt_111 (
    .i_vec(i_mt_l111), .stride(stride_l111), .o_vec(o_mt_l111)
);

// Shifter 112
wire [112*WORD_WIDTH-1:0] i_lifm_l112;
wire [112*WORD_WIDTH-1:0] o_lifm_l112;
wire [112*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l112;
wire [112*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l112;
wire [6:0] stride_l112;

assign i_lifm_l112 = {lifm_line_arr[111], 111*WORD_WIDTH'b0};
assign i_mt_l112 = {mt_line_arr[111], 111*WORD_WIDTH'b0};
assign stride_l112 = psum_arr[111][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(112), .NUMEL_LOG(7)
) vs_lifm_112 (
    .i_vec(i_lifm_l112), .stride(stride_l112), .o_vec(o_lifm_l112)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(112), .NUMEL_LOG(7)
) vs_mt_112 (
    .i_vec(i_mt_l112), .stride(stride_l112), .o_vec(o_mt_l112)
);

// Shifter 113
wire [113*WORD_WIDTH-1:0] i_lifm_l113;
wire [113*WORD_WIDTH-1:0] o_lifm_l113;
wire [113*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l113;
wire [113*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l113;
wire [6:0] stride_l113;

assign i_lifm_l113 = {lifm_line_arr[112], 112*WORD_WIDTH'b0};
assign i_mt_l113 = {mt_line_arr[112], 112*WORD_WIDTH'b0};
assign stride_l113 = psum_arr[112][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(113), .NUMEL_LOG(7)
) vs_lifm_113 (
    .i_vec(i_lifm_l113), .stride(stride_l113), .o_vec(o_lifm_l113)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(113), .NUMEL_LOG(7)
) vs_mt_113 (
    .i_vec(i_mt_l113), .stride(stride_l113), .o_vec(o_mt_l113)
);

// Shifter 114
wire [114*WORD_WIDTH-1:0] i_lifm_l114;
wire [114*WORD_WIDTH-1:0] o_lifm_l114;
wire [114*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l114;
wire [114*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l114;
wire [6:0] stride_l114;

assign i_lifm_l114 = {lifm_line_arr[113], 113*WORD_WIDTH'b0};
assign i_mt_l114 = {mt_line_arr[113], 113*WORD_WIDTH'b0};
assign stride_l114 = psum_arr[113][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(114), .NUMEL_LOG(7)
) vs_lifm_114 (
    .i_vec(i_lifm_l114), .stride(stride_l114), .o_vec(o_lifm_l114)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(114), .NUMEL_LOG(7)
) vs_mt_114 (
    .i_vec(i_mt_l114), .stride(stride_l114), .o_vec(o_mt_l114)
);

// Shifter 115
wire [115*WORD_WIDTH-1:0] i_lifm_l115;
wire [115*WORD_WIDTH-1:0] o_lifm_l115;
wire [115*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l115;
wire [115*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l115;
wire [6:0] stride_l115;

assign i_lifm_l115 = {lifm_line_arr[114], 114*WORD_WIDTH'b0};
assign i_mt_l115 = {mt_line_arr[114], 114*WORD_WIDTH'b0};
assign stride_l115 = psum_arr[114][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(115), .NUMEL_LOG(7)
) vs_lifm_115 (
    .i_vec(i_lifm_l115), .stride(stride_l115), .o_vec(o_lifm_l115)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(115), .NUMEL_LOG(7)
) vs_mt_115 (
    .i_vec(i_mt_l115), .stride(stride_l115), .o_vec(o_mt_l115)
);

// Shifter 116
wire [116*WORD_WIDTH-1:0] i_lifm_l116;
wire [116*WORD_WIDTH-1:0] o_lifm_l116;
wire [116*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l116;
wire [116*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l116;
wire [6:0] stride_l116;

assign i_lifm_l116 = {lifm_line_arr[115], 115*WORD_WIDTH'b0};
assign i_mt_l116 = {mt_line_arr[115], 115*WORD_WIDTH'b0};
assign stride_l116 = psum_arr[115][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(116), .NUMEL_LOG(7)
) vs_lifm_116 (
    .i_vec(i_lifm_l116), .stride(stride_l116), .o_vec(o_lifm_l116)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(116), .NUMEL_LOG(7)
) vs_mt_116 (
    .i_vec(i_mt_l116), .stride(stride_l116), .o_vec(o_mt_l116)
);

// Shifter 117
wire [117*WORD_WIDTH-1:0] i_lifm_l117;
wire [117*WORD_WIDTH-1:0] o_lifm_l117;
wire [117*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l117;
wire [117*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l117;
wire [6:0] stride_l117;

assign i_lifm_l117 = {lifm_line_arr[116], 116*WORD_WIDTH'b0};
assign i_mt_l117 = {mt_line_arr[116], 116*WORD_WIDTH'b0};
assign stride_l117 = psum_arr[116][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(117), .NUMEL_LOG(7)
) vs_lifm_117 (
    .i_vec(i_lifm_l117), .stride(stride_l117), .o_vec(o_lifm_l117)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(117), .NUMEL_LOG(7)
) vs_mt_117 (
    .i_vec(i_mt_l117), .stride(stride_l117), .o_vec(o_mt_l117)
);

// Shifter 118
wire [118*WORD_WIDTH-1:0] i_lifm_l118;
wire [118*WORD_WIDTH-1:0] o_lifm_l118;
wire [118*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l118;
wire [118*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l118;
wire [6:0] stride_l118;

assign i_lifm_l118 = {lifm_line_arr[117], 117*WORD_WIDTH'b0};
assign i_mt_l118 = {mt_line_arr[117], 117*WORD_WIDTH'b0};
assign stride_l118 = psum_arr[117][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(118), .NUMEL_LOG(7)
) vs_lifm_118 (
    .i_vec(i_lifm_l118), .stride(stride_l118), .o_vec(o_lifm_l118)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(118), .NUMEL_LOG(7)
) vs_mt_118 (
    .i_vec(i_mt_l118), .stride(stride_l118), .o_vec(o_mt_l118)
);

// Shifter 119
wire [119*WORD_WIDTH-1:0] i_lifm_l119;
wire [119*WORD_WIDTH-1:0] o_lifm_l119;
wire [119*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l119;
wire [119*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l119;
wire [6:0] stride_l119;

assign i_lifm_l119 = {lifm_line_arr[118], 118*WORD_WIDTH'b0};
assign i_mt_l119 = {mt_line_arr[118], 118*WORD_WIDTH'b0};
assign stride_l119 = psum_arr[118][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(119), .NUMEL_LOG(7)
) vs_lifm_119 (
    .i_vec(i_lifm_l119), .stride(stride_l119), .o_vec(o_lifm_l119)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(119), .NUMEL_LOG(7)
) vs_mt_119 (
    .i_vec(i_mt_l119), .stride(stride_l119), .o_vec(o_mt_l119)
);

// Shifter 120
wire [120*WORD_WIDTH-1:0] i_lifm_l120;
wire [120*WORD_WIDTH-1:0] o_lifm_l120;
wire [120*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l120;
wire [120*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l120;
wire [6:0] stride_l120;

assign i_lifm_l120 = {lifm_line_arr[119], 119*WORD_WIDTH'b0};
assign i_mt_l120 = {mt_line_arr[119], 119*WORD_WIDTH'b0};
assign stride_l120 = psum_arr[119][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(120), .NUMEL_LOG(7)
) vs_lifm_120 (
    .i_vec(i_lifm_l120), .stride(stride_l120), .o_vec(o_lifm_l120)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(120), .NUMEL_LOG(7)
) vs_mt_120 (
    .i_vec(i_mt_l120), .stride(stride_l120), .o_vec(o_mt_l120)
);

// Shifter 121
wire [121*WORD_WIDTH-1:0] i_lifm_l121;
wire [121*WORD_WIDTH-1:0] o_lifm_l121;
wire [121*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l121;
wire [121*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l121;
wire [6:0] stride_l121;

assign i_lifm_l121 = {lifm_line_arr[120], 120*WORD_WIDTH'b0};
assign i_mt_l121 = {mt_line_arr[120], 120*WORD_WIDTH'b0};
assign stride_l121 = psum_arr[120][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(121), .NUMEL_LOG(7)
) vs_lifm_121 (
    .i_vec(i_lifm_l121), .stride(stride_l121), .o_vec(o_lifm_l121)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(121), .NUMEL_LOG(7)
) vs_mt_121 (
    .i_vec(i_mt_l121), .stride(stride_l121), .o_vec(o_mt_l121)
);

// Shifter 122
wire [122*WORD_WIDTH-1:0] i_lifm_l122;
wire [122*WORD_WIDTH-1:0] o_lifm_l122;
wire [122*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l122;
wire [122*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l122;
wire [6:0] stride_l122;

assign i_lifm_l122 = {lifm_line_arr[121], 121*WORD_WIDTH'b0};
assign i_mt_l122 = {mt_line_arr[121], 121*WORD_WIDTH'b0};
assign stride_l122 = psum_arr[121][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(122), .NUMEL_LOG(7)
) vs_lifm_122 (
    .i_vec(i_lifm_l122), .stride(stride_l122), .o_vec(o_lifm_l122)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(122), .NUMEL_LOG(7)
) vs_mt_122 (
    .i_vec(i_mt_l122), .stride(stride_l122), .o_vec(o_mt_l122)
);

// Shifter 123
wire [123*WORD_WIDTH-1:0] i_lifm_l123;
wire [123*WORD_WIDTH-1:0] o_lifm_l123;
wire [123*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l123;
wire [123*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l123;
wire [6:0] stride_l123;

assign i_lifm_l123 = {lifm_line_arr[122], 122*WORD_WIDTH'b0};
assign i_mt_l123 = {mt_line_arr[122], 122*WORD_WIDTH'b0};
assign stride_l123 = psum_arr[122][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(123), .NUMEL_LOG(7)
) vs_lifm_123 (
    .i_vec(i_lifm_l123), .stride(stride_l123), .o_vec(o_lifm_l123)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(123), .NUMEL_LOG(7)
) vs_mt_123 (
    .i_vec(i_mt_l123), .stride(stride_l123), .o_vec(o_mt_l123)
);

// Shifter 124
wire [124*WORD_WIDTH-1:0] i_lifm_l124;
wire [124*WORD_WIDTH-1:0] o_lifm_l124;
wire [124*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l124;
wire [124*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l124;
wire [6:0] stride_l124;

assign i_lifm_l124 = {lifm_line_arr[123], 123*WORD_WIDTH'b0};
assign i_mt_l124 = {mt_line_arr[123], 123*WORD_WIDTH'b0};
assign stride_l124 = psum_arr[123][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(124), .NUMEL_LOG(7)
) vs_lifm_124 (
    .i_vec(i_lifm_l124), .stride(stride_l124), .o_vec(o_lifm_l124)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(124), .NUMEL_LOG(7)
) vs_mt_124 (
    .i_vec(i_mt_l124), .stride(stride_l124), .o_vec(o_mt_l124)
);

// Shifter 125
wire [125*WORD_WIDTH-1:0] i_lifm_l125;
wire [125*WORD_WIDTH-1:0] o_lifm_l125;
wire [125*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l125;
wire [125*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l125;
wire [6:0] stride_l125;

assign i_lifm_l125 = {lifm_line_arr[124], 124*WORD_WIDTH'b0};
assign i_mt_l125 = {mt_line_arr[124], 124*WORD_WIDTH'b0};
assign stride_l125 = psum_arr[124][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(125), .NUMEL_LOG(7)
) vs_lifm_125 (
    .i_vec(i_lifm_l125), .stride(stride_l125), .o_vec(o_lifm_l125)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(125), .NUMEL_LOG(7)
) vs_mt_125 (
    .i_vec(i_mt_l125), .stride(stride_l125), .o_vec(o_mt_l125)
);

// Shifter 126
wire [126*WORD_WIDTH-1:0] i_lifm_l126;
wire [126*WORD_WIDTH-1:0] o_lifm_l126;
wire [126*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l126;
wire [126*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l126;
wire [6:0] stride_l126;

assign i_lifm_l126 = {lifm_line_arr[125], 125*WORD_WIDTH'b0};
assign i_mt_l126 = {mt_line_arr[125], 125*WORD_WIDTH'b0};
assign stride_l126 = psum_arr[125][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(126), .NUMEL_LOG(7)
) vs_lifm_126 (
    .i_vec(i_lifm_l126), .stride(stride_l126), .o_vec(o_lifm_l126)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(126), .NUMEL_LOG(7)
) vs_mt_126 (
    .i_vec(i_mt_l126), .stride(stride_l126), .o_vec(o_mt_l126)
);

// Shifter 127
wire [127*WORD_WIDTH-1:0] i_lifm_l127;
wire [127*WORD_WIDTH-1:0] o_lifm_l127;
wire [127*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l127;
wire [127*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l127;
wire [6:0] stride_l127;

assign i_lifm_l127 = {lifm_line_arr[126], 126*WORD_WIDTH'b0};
assign i_mt_l127 = {mt_line_arr[126], 126*WORD_WIDTH'b0};
assign stride_l127 = psum_arr[126][6:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(127), .NUMEL_LOG(7)
) vs_lifm_127 (
    .i_vec(i_lifm_l127), .stride(stride_l127), .o_vec(o_lifm_l127)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(127), .NUMEL_LOG(7)
) vs_mt_127 (
    .i_vec(i_mt_l127), .stride(stride_l127), .o_vec(o_mt_l127)
);

// Shifter 128
wire [128*WORD_WIDTH-1:0] i_lifm_l128;
wire [128*WORD_WIDTH-1:0] o_lifm_l128;
wire [128*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] i_mt_l128;
wire [128*DIST_WIDTH*MAX_LIFM_RSIZ-1:0] o_mt_l128;
wire [7:0] stride_l128;

assign i_lifm_l128 = {lifm_line_arr[127], 127*WORD_WIDTH'b0};
assign i_mt_l128 = {mt_line_arr[127], 127*WORD_WIDTH'b0};
assign stride_l128 = psum_arr[127][7:0];

VShifter #(
    .WORD_WIDTH(WORD_WIDTH), .NUMEL(128), .NUMEL_LOG(8)
) vs_lifm_128 (
    .i_vec(i_lifm_l128), .stride(stride_l128), .o_vec(o_lifm_l128)
);

VShifter #(
    .WORD_WIDTH(DIST_WIDTH*MAX_LIFM_RSIZ), .NUMEL(128), .NUMEL_LOG(8)
) vs_mt_128 (
    .i_vec(i_mt_l128), .stride(stride_l128), .o_vec(o_mt_l128)
);

assign lifm_comp[0] = o_lifm_l2[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l3[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l4[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l5[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l6[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l7[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l8[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l9[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[0*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[0*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[0]   = o_mt_l2[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l3[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l4[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l5[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l6[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l7[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l8[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l9[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[0*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[1] = o_lifm_l2[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l3[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l4[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l5[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l6[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l7[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l8[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l9[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[1*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[1*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[1]   = o_mt_l2[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l3[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l4[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l5[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l6[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l7[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l8[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l9[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[1*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[2] = o_lifm_l3[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l4[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l5[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l6[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l7[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l8[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l9[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[2*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[2*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[2]   = o_mt_l3[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l4[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l5[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l6[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l7[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l8[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l9[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[2*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[3] = o_lifm_l4[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l5[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l6[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l7[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l8[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l9[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[3*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[3*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[3]   = o_mt_l4[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l5[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l6[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l7[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l8[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l9[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[3*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[4] = o_lifm_l5[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l6[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l7[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l8[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l9[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[4*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[4*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[4]   = o_mt_l5[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l6[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l7[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l8[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l9[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[4*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[5] = o_lifm_l6[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l7[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l8[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l9[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[5*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[5*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[5]   = o_mt_l6[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l7[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l8[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l9[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[5*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[6] = o_lifm_l7[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l8[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l9[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[6*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[6*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[6]   = o_mt_l7[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l8[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l9[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[6*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[7] = o_lifm_l8[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l9[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[7*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[7*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[7]   = o_mt_l8[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l9[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[7*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[8] = o_lifm_l9[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l10[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[8*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[8*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[8]   = o_mt_l9[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l10[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[8*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[9] = o_lifm_l10[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l11[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[9*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[9*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[9]   = o_mt_l10[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l11[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[9*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[10] = o_lifm_l11[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l12[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[10*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[10*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[10]   = o_mt_l11[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l12[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[10*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[11] = o_lifm_l12[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l13[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[11*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[11*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[11]   = o_mt_l12[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l13[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[11*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[12] = o_lifm_l13[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l14[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[12*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[12*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[12]   = o_mt_l13[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l14[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[12*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[13] = o_lifm_l14[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l15[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[13*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[13*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[13]   = o_mt_l14[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l15[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[13*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[14] = o_lifm_l15[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l16[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[14*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[14*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[14]   = o_mt_l15[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l16[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[14*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[15] = o_lifm_l16[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l17[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[15*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[15*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[15]   = o_mt_l16[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l17[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[15*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[16] = o_lifm_l17[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l18[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[16*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[16*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[16]   = o_mt_l17[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l18[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[16*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[17] = o_lifm_l18[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l19[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[17*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[17*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[17]   = o_mt_l18[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l19[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[17*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[18] = o_lifm_l19[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l20[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[18*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[18*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[18]   = o_mt_l19[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l20[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[18*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[19] = o_lifm_l20[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l21[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[19*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[19*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[19]   = o_mt_l20[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l21[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[19*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[20] = o_lifm_l21[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l22[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[20*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[20*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[20]   = o_mt_l21[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l22[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[20*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[21] = o_lifm_l22[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l23[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[21*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[21*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[21]   = o_mt_l22[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l23[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[21*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[22] = o_lifm_l23[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l24[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[22*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[22*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[22]   = o_mt_l23[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l24[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[22*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[23] = o_lifm_l24[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l25[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[23*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[23*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[23]   = o_mt_l24[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l25[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[23*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[24] = o_lifm_l25[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l26[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[24*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[24*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[24]   = o_mt_l25[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l26[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[24*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[25] = o_lifm_l26[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l27[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[25*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[25*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[25]   = o_mt_l26[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l27[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[25*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[26] = o_lifm_l27[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l28[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[26*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[26*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[26]   = o_mt_l27[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l28[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[26*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[27] = o_lifm_l28[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l29[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[27*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[27*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[27]   = o_mt_l28[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l29[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[27*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[28] = o_lifm_l29[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l30[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[28*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[28*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[28]   = o_mt_l29[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l30[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[28*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[29] = o_lifm_l30[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l31[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[29*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[29*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[29]   = o_mt_l30[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l31[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[29*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[30] = o_lifm_l31[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l32[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[30*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[30*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[30]   = o_mt_l31[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l32[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[30*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[31] = o_lifm_l32[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l33[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[31*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[31*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[31]   = o_mt_l32[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l33[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[31*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[32] = o_lifm_l33[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l34[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[32*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[32*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[32]   = o_mt_l33[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l34[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[32*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[33] = o_lifm_l34[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l35[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[33*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[33*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[33]   = o_mt_l34[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l35[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[33*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[34] = o_lifm_l35[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l36[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[34*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[34*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[34]   = o_mt_l35[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l36[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[34*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[35] = o_lifm_l36[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l37[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[35*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[35*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[35]   = o_mt_l36[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l37[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[35*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[36] = o_lifm_l37[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l38[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[36*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[36*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[36]   = o_mt_l37[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l38[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[36*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[37] = o_lifm_l38[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l39[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[37*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[37*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[37]   = o_mt_l38[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l39[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[37*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[38] = o_lifm_l39[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l40[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[38*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[38*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[38]   = o_mt_l39[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l40[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[38*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[39] = o_lifm_l40[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l41[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[39*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[39*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[39]   = o_mt_l40[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l41[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[39*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[40] = o_lifm_l41[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l42[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[40*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[40*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[40]   = o_mt_l41[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l42[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[40*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[41] = o_lifm_l42[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l43[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[41*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[41*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[41]   = o_mt_l42[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l43[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[41*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[42] = o_lifm_l43[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l44[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[42*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[42*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[42]   = o_mt_l43[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l44[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[42*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[43] = o_lifm_l44[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l45[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[43*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[43*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[43]   = o_mt_l44[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l45[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[43*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[44] = o_lifm_l45[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l46[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[44*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[44*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[44]   = o_mt_l45[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l46[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[44*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[45] = o_lifm_l46[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l47[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[45*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[45*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[45]   = o_mt_l46[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l47[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[45*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[46] = o_lifm_l47[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l48[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[46*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[46*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[46]   = o_mt_l47[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l48[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[46*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[47] = o_lifm_l48[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l49[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[47*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[47*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[47]   = o_mt_l48[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l49[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[47*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[48] = o_lifm_l49[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l50[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[48*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[48*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[48]   = o_mt_l49[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l50[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[48*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[49] = o_lifm_l50[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l51[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[49*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[49*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[49]   = o_mt_l50[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l51[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[49*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[50] = o_lifm_l51[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l52[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[50*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[50*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[50]   = o_mt_l51[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l52[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[50*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[51] = o_lifm_l52[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l53[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[51*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[51*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[51]   = o_mt_l52[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l53[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[51*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[52] = o_lifm_l53[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l54[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[52*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[52*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[52]   = o_mt_l53[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l54[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[52*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[53] = o_lifm_l54[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l55[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[53*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[53*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[53]   = o_mt_l54[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l55[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[53*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[54] = o_lifm_l55[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l56[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[54*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[54*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[54]   = o_mt_l55[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l56[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[54*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[55] = o_lifm_l56[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l57[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[55*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[55*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[55]   = o_mt_l56[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l57[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[55*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[56] = o_lifm_l57[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l58[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[56*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[56*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[56]   = o_mt_l57[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l58[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[56*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[57] = o_lifm_l58[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l59[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[57*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[57*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[57]   = o_mt_l58[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l59[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[57*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[58] = o_lifm_l59[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l60[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[58*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[58*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[58]   = o_mt_l59[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l60[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[58*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[59] = o_lifm_l60[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l61[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[59*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[59*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[59]   = o_mt_l60[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l61[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[59*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[60] = o_lifm_l61[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l62[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[60*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[60*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[60]   = o_mt_l61[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l62[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[60*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[61] = o_lifm_l62[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l63[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[61*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[61*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[61]   = o_mt_l62[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l63[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[61*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[62] = o_lifm_l63[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l64[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[62*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[62*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[62]   = o_mt_l63[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l64[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[62*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[63] = o_lifm_l64[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l65[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[63*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[63*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[63]   = o_mt_l64[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l65[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[63*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[64] = o_lifm_l65[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l66[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[64*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[64*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[64]   = o_mt_l65[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l66[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[64*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[65] = o_lifm_l66[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l67[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[65*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[65*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[65]   = o_mt_l66[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l67[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[65*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[66] = o_lifm_l67[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l68[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[66*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[66*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[66]   = o_mt_l67[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l68[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[66*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[67] = o_lifm_l68[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l69[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[67*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[67*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[67]   = o_mt_l68[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l69[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[67*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[68] = o_lifm_l69[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l70[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[68*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[68*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[68]   = o_mt_l69[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l70[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[68*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[69] = o_lifm_l70[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l71[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[69*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[69*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[69]   = o_mt_l70[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l71[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[69*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[70] = o_lifm_l71[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l72[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[70*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[70*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[70]   = o_mt_l71[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l72[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[70*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[71] = o_lifm_l72[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l73[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[71*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[71*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[71]   = o_mt_l72[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l73[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[71*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[72] = o_lifm_l73[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l74[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[72*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[72*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[72]   = o_mt_l73[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l74[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[72*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[73] = o_lifm_l74[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l75[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[73*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[73*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[73]   = o_mt_l74[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l75[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[73*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[74] = o_lifm_l75[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l76[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[74*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[74*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[74]   = o_mt_l75[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l76[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[74*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[75] = o_lifm_l76[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l77[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[75*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[75*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[75]   = o_mt_l76[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l77[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[75*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[76] = o_lifm_l77[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l78[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[76*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[76*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[76]   = o_mt_l77[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l78[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[76*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[77] = o_lifm_l78[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l79[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[77*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[77*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[77]   = o_mt_l78[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l79[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[77*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[78] = o_lifm_l79[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l80[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[78*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[78*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[78]   = o_mt_l79[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l80[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[78*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[79] = o_lifm_l80[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l81[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[79*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[79*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[79]   = o_mt_l80[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l81[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[79*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[80] = o_lifm_l81[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l82[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[80*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[80*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[80]   = o_mt_l81[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l82[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[80*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[81] = o_lifm_l82[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l83[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[81*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[81*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[81]   = o_mt_l82[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l83[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[81*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[82] = o_lifm_l83[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l84[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[82*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[82*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[82]   = o_mt_l83[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l84[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[82*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[83] = o_lifm_l84[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l85[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[83*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[83*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[83]   = o_mt_l84[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l85[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[83*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[84] = o_lifm_l85[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l86[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[84*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[84*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[84]   = o_mt_l85[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l86[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[84*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[85] = o_lifm_l86[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l87[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[85*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[85*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[85]   = o_mt_l86[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l87[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[85*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[86] = o_lifm_l87[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l88[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[86*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[86*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[86]   = o_mt_l87[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l88[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[86*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[87] = o_lifm_l88[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l89[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[87*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[87*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[87]   = o_mt_l88[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l89[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[87*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[88] = o_lifm_l89[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l90[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[88*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[88*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[88]   = o_mt_l89[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l90[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[88*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[89] = o_lifm_l90[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l91[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[89*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[89*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[89]   = o_mt_l90[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l91[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[89*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[90] = o_lifm_l91[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l92[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[90*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[90*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[90]   = o_mt_l91[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l92[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[90*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[91] = o_lifm_l92[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l93[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[91*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[91*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[91]   = o_mt_l92[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l93[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[91*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[92] = o_lifm_l93[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l94[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[92*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[92*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[92]   = o_mt_l93[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l94[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[92*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[93] = o_lifm_l94[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l95[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[93*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[93*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[93]   = o_mt_l94[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l95[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[93*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[94] = o_lifm_l95[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l96[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[94*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[94*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[94]   = o_mt_l95[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l96[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[94*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[95] = o_lifm_l96[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l97[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[95*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[95*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[95]   = o_mt_l96[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l97[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[95*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[96] = o_lifm_l97[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l98[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[96*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[96*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[96]   = o_mt_l97[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l98[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[96*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[97] = o_lifm_l98[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l99[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[97*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[97*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[97]   = o_mt_l98[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l99[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[97*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[98] = o_lifm_l99[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l100[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[98*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[98*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[98]   = o_mt_l99[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l100[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[98*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[99] = o_lifm_l100[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l101[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[99*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[99*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[99]   = o_mt_l100[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l101[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[99*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[100] = o_lifm_l101[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l102[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[100*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[100*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[100]   = o_mt_l101[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l102[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[100*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[101] = o_lifm_l102[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l103[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[101*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[101*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[101]   = o_mt_l102[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l103[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[101*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[102] = o_lifm_l103[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l104[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[102*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[102*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[102]   = o_mt_l103[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l104[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[102*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[103] = o_lifm_l104[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l105[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[103*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[103*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[103]   = o_mt_l104[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l105[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[103*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[104] = o_lifm_l105[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l106[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[104*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[104*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[104]   = o_mt_l105[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l106[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[104*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[105] = o_lifm_l106[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l107[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[105*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[105*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[105]   = o_mt_l106[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l107[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[105*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[106] = o_lifm_l107[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l108[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[106*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[106*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[106]   = o_mt_l107[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l108[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[106*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[107] = o_lifm_l108[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l109[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[107*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[107*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[107]   = o_mt_l108[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l109[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[107*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[108] = o_lifm_l109[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l110[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[108*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[108*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[108]   = o_mt_l109[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l110[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[108*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[109] = o_lifm_l110[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l111[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[109*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[109*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[109]   = o_mt_l110[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l111[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[109*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[110] = o_lifm_l111[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l112[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[110*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[110*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[110]   = o_mt_l111[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l112[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[110*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[111] = o_lifm_l112[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l113[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[111*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[111*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[111]   = o_mt_l112[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l113[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[111*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[112] = o_lifm_l113[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l114[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[112*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[112*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[112]   = o_mt_l113[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l114[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[112*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[113] = o_lifm_l114[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l115[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[113*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[113*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[113]   = o_mt_l114[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l115[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[113*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[114] = o_lifm_l115[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l116[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[114*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[114*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[114]   = o_mt_l115[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l116[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[114*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[115] = o_lifm_l116[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l117[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[115*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[115*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[115]   = o_mt_l116[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l117[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[115*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[116] = o_lifm_l117[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l118[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[116*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[116*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[116]   = o_mt_l117[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l118[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[116*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[117] = o_lifm_l118[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l119[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[117*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[117*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[117]   = o_mt_l118[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l119[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[117*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[118] = o_lifm_l119[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l120[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[118*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[118*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[118]   = o_mt_l119[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l120[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[118*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[119] = o_lifm_l120[119*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l121[119*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[119*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[119*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[119*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[119*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[119*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[119*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[119*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[119]   = o_mt_l120[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l121[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[119*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[120] = o_lifm_l121[120*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l122[120*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[120*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[120*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[120*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[120*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[120*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[120*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[120]   = o_mt_l121[120*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l122[120*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[120*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[120*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[120*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[120*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[120*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[120*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[121] = o_lifm_l122[121*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l123[121*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[121*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[121*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[121*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[121*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[121*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[121]   = o_mt_l122[121*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l123[121*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[121*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[121*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[121*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[121*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[121*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[122] = o_lifm_l123[122*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l124[122*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[122*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[122*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[122*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[122*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[122]   = o_mt_l123[122*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l124[122*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[122*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[122*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[122*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[122*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[123] = o_lifm_l124[123*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l125[123*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[123*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[123*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[123*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[123]   = o_mt_l124[123*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l125[123*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[123*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[123*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[123*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[124] = o_lifm_l125[124*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l126[124*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[124*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[124*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[124]   = o_mt_l125[124*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l126[124*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[124*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[124*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[125] = o_lifm_l126[125*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l127[125*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[125*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[125]   = o_mt_l126[125*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l127[125*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[125*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[126] = o_lifm_l127[126*WORD_WIDTH+:WORD_WIDTH] | o_lifm_l128[126*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[126]   = o_mt_l127[126*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ] | o_mt_l128[126*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]
assign lifm_comp[127] = o_lifm_l128[127*WORD_WIDTH+:WORD_WIDTH]
assign mt_comp[127]   = o_mt_l128[127*DIST_WIDTH*MAX_LIFM_RSIZ+:DIST_WIDTH*MAX_LIFM_RSIZ]

endmodule


module VShifter #(
    parameter WORD_WIDTH = 8,
    parameter NUMEL      = 128,
    parameter NUMEL_LOG  = 7
) (
    input [WORD_WIDTH*NUMEL-1:0] i_vec,
    input [NUMEL_LOG-1:0]        stride,

    output [WORD_WIDTH*NUMEL-1:0] o_vec
);

assign o_vec = i_vec >> (stride * WORD_WIDTH);
    
endmodule